module bondpad_70x70 (
  inout pad
);

endmodule