module neorv32_cpu_cp_muldiv_3f29546453678b855931c174a97d6c0894b8f546
  (input  clk_i,
   input  rstn_i,
   input  \ctrl_i_ctrl_i[if_fence] ,
   input  \ctrl_i_ctrl_i[rf_wb_en] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs1] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs2] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rd] ,
   input  \ctrl_i_ctrl_i[rf_zero_we] ,
   input  [2:0] \ctrl_i_ctrl_i[alu_op] ,
   input  \ctrl_i_ctrl_i[alu_sub] ,
   input  \ctrl_i_ctrl_i[alu_opa_mux] ,
   input  \ctrl_i_ctrl_i[alu_opb_mux] ,
   input  \ctrl_i_ctrl_i[alu_unsigned] ,
   input  \ctrl_i_ctrl_i[alu_cp_alu] ,
   input  \ctrl_i_ctrl_i[alu_cp_cfu] ,
   input  \ctrl_i_ctrl_i[alu_cp_fpu] ,
   input  \ctrl_i_ctrl_i[lsu_req] ,
   input  \ctrl_i_ctrl_i[lsu_rw] ,
   input  \ctrl_i_ctrl_i[lsu_mo_we] ,
   input  \ctrl_i_ctrl_i[lsu_fence] ,
   input  \ctrl_i_ctrl_i[lsu_priv] ,
   input  [2:0] \ctrl_i_ctrl_i[ir_funct3] ,
   input  [11:0] \ctrl_i_ctrl_i[ir_funct12] ,
   input  [6:0] \ctrl_i_ctrl_i[ir_opcode] ,
   input  \ctrl_i_ctrl_i[cpu_priv] ,
   input  \ctrl_i_ctrl_i[cpu_sleep] ,
   input  \ctrl_i_ctrl_i[cpu_trap] ,
   input  \ctrl_i_ctrl_i[cpu_debug] ,
   input  [31:0] rs1_i,
   input  [31:0] rs2_i,
   output [31:0] res_o,
   output valid_o);
  wire [58:0] n15221;
  wire valid_cmd;
  wire [9:0] ctrl;
  wire [194:0] div;
  wire [230:0] mul;
  wire n15225;
  wire n15226;
  wire n15227;
  wire [6:0] n15228;
  wire n15230;
  wire n15231;
  wire n15232;
  wire n15233;
  wire n15234;
  wire n15236;
  wire n15237;
  wire n15238;
  wire n15239;
  wire n15242;
  wire [1:0] n15249;
  wire [1:0] n15253;
  wire [1:0] n15254;
  wire n15256;
  wire [4:0] n15257;
  wire [4:0] n15259;
  wire n15267;
  wire n15269;
  wire n15271;
  wire n15272;
  wire n15273;
  wire n15274;
  wire n15275;
  wire n15276;
  wire n15277;
  wire n15278;
  wire n15279;
  wire n15280;
  wire n15281;
  wire [1:0] n15283;
  wire [1:0] n15284;
  wire n15286;
  wire [1:0] n15289;
  reg [1:0] n15290;
  reg [4:0] n15291;
  reg n15292;
  wire [6:0] n15293;
  wire [6:0] n15298;
  wire [1:0] n15303;
  wire n15305;
  wire n15306;
  wire [2:0] n15309;
  wire n15311;
  wire [2:0] n15312;
  wire n15314;
  wire n15315;
  wire [2:0] n15316;
  wire n15318;
  wire n15319;
  wire [2:0] n15320;
  wire n15322;
  wire n15323;
  wire n15324;
  wire [2:0] n15327;
  wire n15329;
  wire [2:0] n15330;
  wire n15332;
  wire n15333;
  wire [2:0] n15334;
  wire n15336;
  wire n15337;
  wire n15338;
  wire n15341;
  wire n15342;
  wire n15343;
  wire n15344;
  wire n15347;
  wire n15348;
  wire n15349;
  wire n15355;
  wire n15358;
  wire [1:0] n15360;
  wire n15362;
  wire [32:0] n15363;
  wire [30:0] n15364;
  wire [63:0] n15365;
  wire [63:0] n15366;
  wire [63:0] n15367;
  wire [63:0] n15368;
  wire [63:0] n15369;
  wire n15375;
  wire [1:0] n15376;
  wire n15378;
  wire n15379;
  wire n15380;
  wire n15381;
  wire [31:0] n15382;
  wire [32:0] n15383;
  wire n15384;
  wire n15385;
  wire n15386;
  wire [32:0] n15387;
  wire [32:0] n15388;
  wire n15389;
  wire [31:0] n15390;
  wire [32:0] n15391;
  wire n15392;
  wire n15393;
  wire n15394;
  wire [32:0] n15395;
  wire [32:0] n15396;
  wire [32:0] n15397;
  wire n15398;
  wire [31:0] n15399;
  wire [32:0] n15400;
  wire [32:0] n15401;
  wire n15403;
  wire n15404;
  wire n15405;
  wire n15407;
  wire n15413;
  wire n15414;
  wire n15415;
  wire n15416;
  wire [31:0] n15418;
  wire [31:0] n15419;
  wire n15420;
  wire n15421;
  wire n15422;
  wire [31:0] n15424;
  wire [31:0] n15425;
  wire [1:0] n15426;
  wire n15428;
  wire n15429;
  wire n15430;
  wire n15431;
  wire n15438;
  wire n15440;
  wire n15442;
  wire n15443;
  wire n15444;
  wire n15445;
  wire n15446;
  wire n15447;
  wire n15448;
  wire n15449;
  wire n15450;
  wire n15451;
  wire n15452;
  wire n15453;
  wire n15454;
  wire n15455;
  wire n15456;
  wire n15457;
  wire n15458;
  wire n15459;
  wire n15460;
  wire n15461;
  wire n15462;
  wire n15463;
  wire n15464;
  wire n15465;
  wire n15466;
  wire n15467;
  wire n15468;
  wire n15469;
  wire n15470;
  wire n15471;
  wire n15472;
  wire n15473;
  wire n15474;
  wire n15475;
  wire n15476;
  wire n15477;
  wire n15478;
  wire n15479;
  wire n15480;
  wire n15481;
  wire n15482;
  wire n15483;
  wire n15484;
  wire n15485;
  wire n15486;
  wire n15487;
  wire n15488;
  wire n15489;
  wire n15490;
  wire n15491;
  wire n15492;
  wire n15493;
  wire n15494;
  wire n15495;
  wire n15496;
  wire n15497;
  wire n15498;
  wire n15499;
  wire n15500;
  wire n15501;
  wire n15502;
  wire n15503;
  wire n15504;
  wire [1:0] n15505;
  wire n15507;
  wire n15508;
  wire n15510;
  wire n15511;
  wire [1:0] n15513;
  wire n15515;
  wire [1:0] n15516;
  wire n15518;
  wire n15519;
  wire [30:0] n15520;
  wire n15521;
  wire n15522;
  wire [31:0] n15523;
  wire n15524;
  wire n15525;
  wire [31:0] n15526;
  wire [30:0] n15527;
  wire n15528;
  wire [31:0] n15529;
  wire [31:0] n15530;
  wire [63:0] n15531;
  wire [63:0] n15532;
  wire [63:0] n15533;
  wire [96:0] n15534;
  wire [32:0] n15535;
  wire [32:0] n15536;
  wire [32:0] n15537;
  wire [63:0] n15538;
  wire [63:0] n15539;
  wire [96:0] n15540;
  wire [96:0] n15543;
  wire [30:0] n15546;
  wire [31:0] n15548;
  wire n15549;
  wire [32:0] n15550;
  wire [31:0] n15551;
  wire [32:0] n15553;
  wire [32:0] n15554;
  wire [31:0] n15555;
  wire [1:0] n15556;
  wire n15558;
  wire [31:0] n15559;
  wire [31:0] n15560;
  wire [31:0] n15561;
  wire [31:0] n15563;
  wire n15564;
  wire [31:0] n15565;
  wire [31:0] n15566;
  wire n15568;
  wire [2:0] n15569;
  wire [31:0] n15570;
  wire n15572;
  wire [31:0] n15573;
  wire n15575;
  wire n15577;
  wire n15578;
  wire n15580;
  wire n15581;
  wire [31:0] n15582;
  wire [1:0] n15583;
  reg [31:0] n15584;
  wire [31:0] n15586;
  reg n15589;
  reg [6:0] n15590;
  wire [9:0] n15591;
  reg [96:0] n15592;
  wire [194:0] n15593;
  reg [63:0] n15594;
  wire [230:0] n15595;
  assign res_o = n15586; //(module output)
  assign valid_o = n15306; //(module output)
  assign n15221 = {\ctrl_i_ctrl_i[cpu_debug] , \ctrl_i_ctrl_i[cpu_trap] , \ctrl_i_ctrl_i[cpu_sleep] , \ctrl_i_ctrl_i[cpu_priv] , \ctrl_i_ctrl_i[ir_opcode] , \ctrl_i_ctrl_i[ir_funct12] , \ctrl_i_ctrl_i[ir_funct3] , \ctrl_i_ctrl_i[lsu_priv] , \ctrl_i_ctrl_i[lsu_fence] , \ctrl_i_ctrl_i[lsu_mo_we] , \ctrl_i_ctrl_i[lsu_rw] , \ctrl_i_ctrl_i[lsu_req] , \ctrl_i_ctrl_i[alu_cp_fpu] , \ctrl_i_ctrl_i[alu_cp_cfu] , \ctrl_i_ctrl_i[alu_cp_alu] , \ctrl_i_ctrl_i[alu_unsigned] , \ctrl_i_ctrl_i[alu_opb_mux] , \ctrl_i_ctrl_i[alu_opa_mux] , \ctrl_i_ctrl_i[alu_sub] , \ctrl_i_ctrl_i[alu_op] , \ctrl_i_ctrl_i[rf_zero_we] , \ctrl_i_ctrl_i[rf_rd] , \ctrl_i_ctrl_i[rf_rs2] , \ctrl_i_ctrl_i[rf_rs1] , \ctrl_i_ctrl_i[rf_wb_en] , \ctrl_i_ctrl_i[if_fence] };
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:55:10  */
  assign valid_cmd = n15239; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:66:10  */
  assign ctrl = n15591; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:79:10  */
  assign div = n15593; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:91:10  */
  assign mul = n15595; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:97:33  */
  assign n15225 = n15221[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:97:72  */
  assign n15226 = n15221[53]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:97:51  */
  assign n15227 = n15226 & n15225;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:98:43  */
  assign n15228 = n15221[47:41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:98:57  */
  assign n15230 = n15228 == 7'b0000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:97:83  */
  assign n15231 = n15230 & n15227;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:99:43  */
  assign n15232 = n15221[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:99:47  */
  assign n15233 = ~n15232;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:99:75  */
  assign n15234 = n15221[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:99:86  */
  assign n15236 = 1'b1 & n15234;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:99:54  */
  assign n15237 = n15233 | n15236;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:98:70  */
  assign n15238 = n15237 & n15231;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:97:20  */
  assign n15239 = n15238 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:106:16  */
  assign n15242 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:116:17  */
  assign n15249 = ctrl[1:0]; // extract
  assign n15253 = ctrl[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:120:11  */
  assign n15254 = valid_cmd ? 2'b01 : n15253;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:118:9  */
  assign n15256 = n15249 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:130:55  */
  assign n15257 = ctrl[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:130:60  */
  assign n15259 = n15257 - 5'b00001;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15267 = ctrl[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15269 = 1'b0 | n15267;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15271 = ctrl[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15272 = n15269 | n15271;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15273 = ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15274 = n15272 | n15273;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15275 = ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15276 = n15274 | n15275;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15277 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15278 = n15276 | n15277;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:131:37  */
  assign n15279 = ~n15278;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:131:55  */
  assign n15280 = n15221[57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:131:44  */
  assign n15281 = n15279 | n15280;
  assign n15283 = ctrl[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:131:11  */
  assign n15284 = n15281 ? 2'b10 : n15283;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:128:9  */
  assign n15286 = n15249 == 2'b01;
  assign n15289 = {n15286, n15256};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:116:7  */
  always @*
    case (n15289)
      2'b10: n15290 = n15284;
      2'b01: n15290 = n15254;
      default: n15290 = 2'b00;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:116:7  */
  always @*
    case (n15289)
      2'b10: n15291 = n15259;
      2'b01: n15291 = 5'b11110;
      default: n15291 = 5'b11110;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:116:7  */
  always @*
    case (n15289)
      2'b10: n15292 = 1'b0;
      2'b01: n15292 = 1'b0;
      default: n15292 = 1'b1;
    endcase
  assign n15293 = {n15291, n15290};
  assign n15298 = {5'b00000, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:145:29  */
  assign n15303 = ctrl[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:145:35  */
  assign n15305 = n15303 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:145:18  */
  assign n15306 = n15305 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:148:42  */
  assign n15309 = n15221[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:148:52  */
  assign n15311 = n15309 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:148:76  */
  assign n15312 = n15221[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:148:86  */
  assign n15314 = n15312 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:148:65  */
  assign n15315 = n15311 | n15314;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:149:42  */
  assign n15316 = n15221[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:149:52  */
  assign n15318 = n15316 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:148:101  */
  assign n15319 = n15315 | n15318;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:149:76  */
  assign n15320 = n15221[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:149:86  */
  assign n15322 = n15320 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:149:65  */
  assign n15323 = n15319 | n15322;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:148:29  */
  assign n15324 = n15323 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:150:42  */
  assign n15327 = n15221[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:150:52  */
  assign n15329 = n15327 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:151:42  */
  assign n15330 = n15221[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:151:52  */
  assign n15332 = n15330 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:150:65  */
  assign n15333 = n15329 | n15332;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:151:76  */
  assign n15334 = n15221[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:151:86  */
  assign n15336 = n15334 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:151:65  */
  assign n15337 = n15333 | n15336;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:150:29  */
  assign n15338 = n15337 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:154:64  */
  assign n15341 = n15221[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:154:68  */
  assign n15342 = ~n15341;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:154:43  */
  assign n15343 = n15342 & valid_cmd;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:154:20  */
  assign n15344 = n15343 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:155:64  */
  assign n15347 = n15221[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:155:43  */
  assign n15348 = n15347 & valid_cmd;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:155:20  */
  assign n15349 = n15348 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:207:18  */
  assign n15355 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:210:17  */
  assign n15358 = mul[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:213:21  */
  assign n15360 = ctrl[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:213:27  */
  assign n15362 = n15360 != 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:214:44  */
  assign n15363 = mul[97:65]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:215:45  */
  assign n15364 = mul[32:2]; // extract
  assign n15365 = {n15363, n15364};
  assign n15366 = mul[64:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:213:9  */
  assign n15367 = n15362 ? n15365 : n15366;
  assign n15368 = {32'b00000000000000000000000000000000, rs1_i};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:210:9  */
  assign n15369 = n15358 ? n15368 : n15367;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:223:19  */
  assign n15375 = mul[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:224:18  */
  assign n15376 = ctrl[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:224:24  */
  assign n15378 = n15376 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:224:44  */
  assign n15379 = ctrl[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:224:34  */
  assign n15380 = n15379 & n15378;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:225:53  */
  assign n15381 = mul[98]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:225:70  */
  assign n15382 = mul[64:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:225:60  */
  assign n15383 = {n15381, n15382};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:225:103  */
  assign n15384 = rs2_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:225:125  */
  assign n15385 = ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:225:116  */
  assign n15386 = n15384 & n15385;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:225:140  */
  assign n15387 = {n15386, rs2_i};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:225:86  */
  assign n15388 = n15383 - n15387;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:227:53  */
  assign n15389 = mul[98]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:227:70  */
  assign n15390 = mul[64:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:227:60  */
  assign n15391 = {n15389, n15390};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:227:103  */
  assign n15392 = rs2_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:227:125  */
  assign n15393 = ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:227:116  */
  assign n15394 = n15392 & n15393;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:227:140  */
  assign n15395 = {n15394, rs2_i};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:227:86  */
  assign n15396 = n15391 + n15395;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:224:9  */
  assign n15397 = n15380 ? n15388 : n15396;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:230:24  */
  assign n15398 = mul[98]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:230:41  */
  assign n15399 = mul[64:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:230:31  */
  assign n15400 = {n15398, n15399};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:223:7  */
  assign n15401 = n15375 ? n15397 : n15400;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:235:27  */
  assign n15403 = mul[64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:235:52  */
  assign n15404 = ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:235:43  */
  assign n15405 = n15403 & n15404;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:255:18  */
  assign n15407 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:261:17  */
  assign n15413 = div[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:263:21  */
  assign n15414 = rs1_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:263:43  */
  assign n15415 = ctrl[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:263:34  */
  assign n15416 = n15414 & n15415;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:264:49  */
  assign n15418 = 32'b00000000000000000000000000000000 - rs1_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:263:11  */
  assign n15419 = n15416 ? n15418 : rs1_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:269:21  */
  assign n15420 = rs2_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:269:43  */
  assign n15421 = ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:269:34  */
  assign n15422 = n15420 & n15421;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:270:48  */
  assign n15424 = 32'b00000000000000000000000000000000 - rs2_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:269:11  */
  assign n15425 = n15422 ? n15424 : rs2_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:275:31  */
  assign n15426 = n15221[34:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:275:44  */
  assign n15428 = n15426 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:276:35  */
  assign n15429 = rs1_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:276:57  */
  assign n15430 = rs2_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:276:48  */
  assign n15431 = n15429 ^ n15430;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15438 = rs2_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15440 = 1'b0 | n15438;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15442 = rs2_i[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15443 = n15440 | n15442;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15444 = rs2_i[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15445 = n15443 | n15444;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15446 = rs2_i[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15447 = n15445 | n15446;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15448 = rs2_i[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15449 = n15447 | n15448;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15450 = rs2_i[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15451 = n15449 | n15450;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15452 = rs2_i[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15453 = n15451 | n15452;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15454 = rs2_i[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15455 = n15453 | n15454;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15456 = rs2_i[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15457 = n15455 | n15456;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15458 = rs2_i[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15459 = n15457 | n15458;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15460 = rs2_i[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15461 = n15459 | n15460;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15462 = rs2_i[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15463 = n15461 | n15462;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15464 = rs2_i[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15465 = n15463 | n15464;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15466 = rs2_i[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15467 = n15465 | n15466;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15468 = rs2_i[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15469 = n15467 | n15468;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15470 = rs2_i[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15471 = n15469 | n15470;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15472 = rs2_i[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15473 = n15471 | n15472;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15474 = rs2_i[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15475 = n15473 | n15474;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15476 = rs2_i[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15477 = n15475 | n15476;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15478 = rs2_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15479 = n15477 | n15478;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15480 = rs2_i[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15481 = n15479 | n15480;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15482 = rs2_i[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15483 = n15481 | n15482;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15484 = rs2_i[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15485 = n15483 | n15484;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15486 = rs2_i[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15487 = n15485 | n15486;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15488 = rs2_i[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15489 = n15487 | n15488;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15490 = rs2_i[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15491 = n15489 | n15490;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15492 = rs2_i[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15493 = n15491 | n15492;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15494 = rs2_i[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15495 = n15493 | n15494;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15496 = rs2_i[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15497 = n15495 | n15496;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15498 = rs2_i[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15499 = n15497 | n15498;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15500 = rs2_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15501 = n15499 | n15500;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15502 = rs2_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15503 = n15501 | n15502;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:276:71  */
  assign n15504 = n15431 & n15503;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:277:34  */
  assign n15505 = n15221[34:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:277:47  */
  assign n15507 = n15505 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:278:34  */
  assign n15508 = rs1_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:277:11  */
  assign n15510 = n15507 ? n15508 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:275:11  */
  assign n15511 = n15428 ? n15504 : n15510;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:284:21  */
  assign n15513 = ctrl[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:284:27  */
  assign n15515 = n15513 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:284:46  */
  assign n15516 = ctrl[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:284:52  */
  assign n15518 = n15516 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:284:37  */
  assign n15519 = n15515 | n15518;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:285:39  */
  assign n15520 = div[96:66]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:285:67  */
  assign n15521 = div[130]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:285:56  */
  assign n15522 = ~n15521;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:285:53  */
  assign n15523 = {n15520, n15522};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:286:22  */
  assign n15524 = div[130]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:286:27  */
  assign n15525 = ~n15524;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:287:37  */
  assign n15526 = div[129:98]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:289:43  */
  assign n15527 = div[64:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:289:71  */
  assign n15528 = div[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:289:57  */
  assign n15529 = {n15527, n15528};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:286:11  */
  assign n15530 = n15525 ? n15526 : n15529;
  assign n15531 = {n15523, n15530};
  assign n15532 = div[97:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:284:9  */
  assign n15533 = n15519 ? n15531 : n15532;
  assign n15534 = {n15419, 32'b00000000000000000000000000000000, n15425, n15511};
  assign n15535 = n15534[32:0]; // extract
  assign n15536 = div[33:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:261:9  */
  assign n15537 = n15413 ? n15535 : n15536;
  assign n15538 = n15534[96:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:261:9  */
  assign n15539 = n15413 ? n15538 : n15533;
  assign n15540 = {n15539, n15537};
  assign n15543 = {32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:62  */
  assign n15546 = div[64:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:47  */
  assign n15548 = {1'b0, n15546};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:90  */
  assign n15549 = div[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:76  */
  assign n15550 = {n15548, n15549};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:117  */
  assign n15551 = div[33:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:111  */
  assign n15553 = {1'b0, n15551};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:296:96  */
  assign n15554 = n15550 - n15553;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:299:22  */
  assign n15555 = div[97:66]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:299:53  */
  assign n15556 = n15221[35:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:299:66  */
  assign n15558 = n15556 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:299:31  */
  assign n15559 = n15558 ? n15555 : n15560;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:299:99  */
  assign n15560 = div[65:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:300:53  */
  assign n15561 = div[162:131]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:300:38  */
  assign n15563 = 32'b00000000000000000000000000000000 - n15561;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:300:71  */
  assign n15564 = div[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:300:61  */
  assign n15565 = n15564 ? n15563 : n15566;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:300:96  */
  assign n15566 = div[162:131]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:322:14  */
  assign n15568 = ctrl[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:323:19  */
  assign n15569 = n15221[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:325:28  */
  assign n15570 = mul[32:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:324:9  */
  assign n15572 = n15569 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:327:28  */
  assign n15573 = mul[64:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:326:9  */
  assign n15575 = n15569 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:326:24  */
  assign n15577 = n15569 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:326:24  */
  assign n15578 = n15575 | n15577;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:326:38  */
  assign n15580 = n15569 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:326:38  */
  assign n15581 = n15578 | n15580;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:329:24  */
  assign n15582 = div[194:163]; // extract
  assign n15583 = {n15581, n15572};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:323:7  */
  always @*
    case (n15583)
      2'b10: n15584 = n15573;
      2'b01: n15584 = n15570;
      default: n15584 = n15582;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:322:5  */
  assign n15586 = n15568 ? n15584 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:110:5  */
  always @(posedge clk_i or posedge n15242)
    if (n15242)
      n15589 <= 1'b0;
    else
      n15589 <= n15292;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:110:5  */
  always @(posedge clk_i or posedge n15242)
    if (n15242)
      n15590 <= n15298;
    else
      n15590 <= n15293;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:106:5  */
  assign n15591 = {n15589, n15338, n15324, n15590};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:260:7  */
  always @(posedge clk_i or posedge n15407)
    if (n15407)
      n15592 <= n15543;
    else
      n15592 <= n15540;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:255:7  */
  assign n15593 = {n15565, n15559, n15554, n15592, n15349};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:209:7  */
  always @(posedge clk_i or posedge n15355)
    if (n15355)
      n15594 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n15594 <= n15369;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_muldiv.vhd:207:7  */
  assign n15595 = {66'b000000000000000000000000000000000000000000000000000000000000000000, 33'b000000000000000000000000000000000, 33'b000000000000000000000000000000000, n15405, n15401, n15594, n15344};
endmodule

module neorv32_cpu_cp_shifter_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk_i,
   input  rstn_i,
   input  \ctrl_i_ctrl_i[if_fence] ,
   input  \ctrl_i_ctrl_i[rf_wb_en] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs1] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs2] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rd] ,
   input  \ctrl_i_ctrl_i[rf_zero_we] ,
   input  [2:0] \ctrl_i_ctrl_i[alu_op] ,
   input  \ctrl_i_ctrl_i[alu_sub] ,
   input  \ctrl_i_ctrl_i[alu_opa_mux] ,
   input  \ctrl_i_ctrl_i[alu_opb_mux] ,
   input  \ctrl_i_ctrl_i[alu_unsigned] ,
   input  \ctrl_i_ctrl_i[alu_cp_alu] ,
   input  \ctrl_i_ctrl_i[alu_cp_cfu] ,
   input  \ctrl_i_ctrl_i[alu_cp_fpu] ,
   input  \ctrl_i_ctrl_i[lsu_req] ,
   input  \ctrl_i_ctrl_i[lsu_rw] ,
   input  \ctrl_i_ctrl_i[lsu_mo_we] ,
   input  \ctrl_i_ctrl_i[lsu_fence] ,
   input  \ctrl_i_ctrl_i[lsu_priv] ,
   input  [2:0] \ctrl_i_ctrl_i[ir_funct3] ,
   input  [11:0] \ctrl_i_ctrl_i[ir_funct12] ,
   input  [6:0] \ctrl_i_ctrl_i[ir_opcode] ,
   input  \ctrl_i_ctrl_i[cpu_priv] ,
   input  \ctrl_i_ctrl_i[cpu_sleep] ,
   input  \ctrl_i_ctrl_i[cpu_trap] ,
   input  \ctrl_i_ctrl_i[cpu_debug] ,
   input  [31:0] rs1_i,
   input  [4:0] shamt_i,
   output [31:0] res_o,
   output valid_o);
  wire [58:0] n15093;
  wire valid_cmd;
  wire [40:0] shifter;
  wire n15097;
  wire [2:0] n15098;
  wire n15100;
  wire [6:0] n15101;
  wire n15103;
  wire n15104;
  wire [2:0] n15105;
  wire n15107;
  wire [6:0] n15108;
  wire n15110;
  wire n15111;
  wire n15112;
  wire [2:0] n15113;
  wire n15115;
  wire [6:0] n15116;
  wire n15118;
  wire n15119;
  wire n15120;
  wire n15121;
  wire n15122;
  wire n15125;
  wire n15131;
  wire n15132;
  wire n15133;
  wire n15135;
  wire n15136;
  wire n15137;
  wire n15139;
  wire n15140;
  wire n15141;
  wire n15142;
  wire [4:0] n15143;
  wire [4:0] n15145;
  wire n15146;
  wire n15147;
  wire [30:0] n15148;
  wire [31:0] n15150;
  wire n15151;
  wire n15152;
  wire n15153;
  wire [30:0] n15154;
  wire [31:0] n15155;
  wire [31:0] n15156;
  wire [36:0] n15157;
  wire [36:0] n15158;
  wire [36:0] n15159;
  wire [36:0] n15160;
  wire [36:0] n15161;
  wire [37:0] n15162;
  wire [37:0] n15167;
  wire n15178;
  wire n15180;
  wire n15182;
  wire n15183;
  wire n15184;
  wire n15185;
  wire n15186;
  wire n15187;
  wire n15188;
  wire n15189;
  wire n15197;
  wire n15199;
  wire n15201;
  wire n15202;
  wire n15203;
  wire n15204;
  wire n15205;
  wire n15206;
  wire n15207;
  wire n15208;
  wire n15209;
  wire n15210;
  wire [31:0] n15211;
  wire n15212;
  wire [31:0] n15213;
  reg [37:0] n15215;
  reg n15216;
  wire [40:0] n15217;
  assign res_o = n15213; //(module output)
  assign valid_o = n15210; //(module output)
  assign n15093 = {\ctrl_i_ctrl_i[cpu_debug] , \ctrl_i_ctrl_i[cpu_trap] , \ctrl_i_ctrl_i[cpu_sleep] , \ctrl_i_ctrl_i[cpu_priv] , \ctrl_i_ctrl_i[ir_opcode] , \ctrl_i_ctrl_i[ir_funct12] , \ctrl_i_ctrl_i[ir_funct3] , \ctrl_i_ctrl_i[lsu_priv] , \ctrl_i_ctrl_i[lsu_fence] , \ctrl_i_ctrl_i[lsu_mo_we] , \ctrl_i_ctrl_i[lsu_rw] , \ctrl_i_ctrl_i[lsu_req] , \ctrl_i_ctrl_i[alu_cp_fpu] , \ctrl_i_ctrl_i[alu_cp_cfu] , \ctrl_i_ctrl_i[alu_cp_alu] , \ctrl_i_ctrl_i[alu_unsigned] , \ctrl_i_ctrl_i[alu_opb_mux] , \ctrl_i_ctrl_i[alu_opa_mux] , \ctrl_i_ctrl_i[alu_sub] , \ctrl_i_ctrl_i[alu_op] , \ctrl_i_ctrl_i[rf_zero_we] , \ctrl_i_ctrl_i[rf_rd] , \ctrl_i_ctrl_i[rf_rs2] , \ctrl_i_ctrl_i[rf_rs1] , \ctrl_i_ctrl_i[rf_wb_en] , \ctrl_i_ctrl_i[if_fence] };
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:42:10  */
  assign valid_cmd = n15122; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:53:10  */
  assign shifter = n15217; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:65:33  */
  assign n15097 = n15093[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:66:35  */
  assign n15098 = n15093[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:66:45  */
  assign n15100 = n15098 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:66:83  */
  assign n15101 = n15093[47:41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:66:97  */
  assign n15103 = n15101 == 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:66:61  */
  assign n15104 = n15103 & n15100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:67:35  */
  assign n15105 = n15093[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:67:45  */
  assign n15107 = n15105 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:67:83  */
  assign n15108 = n15093[47:41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:67:97  */
  assign n15110 = n15108 == 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:67:61  */
  assign n15111 = n15110 & n15107;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:66:111  */
  assign n15112 = n15104 | n15111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:68:35  */
  assign n15113 = n15093[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:68:45  */
  assign n15115 = n15113 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:68:83  */
  assign n15116 = n15093[47:41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:68:97  */
  assign n15118 = n15116 == 7'b0100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:68:61  */
  assign n15119 = n15118 & n15115;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:67:111  */
  assign n15120 = n15112 | n15119;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:65:51  */
  assign n15121 = n15120 & n15097;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:65:20  */
  assign n15122 = n15121 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:79:18  */
  assign n15125 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:86:36  */
  assign n15131 = shifter[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:86:53  */
  assign n15132 = shifter[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:86:41  */
  assign n15133 = n15131 & n15132;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:89:24  */
  assign n15135 = shifter[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:89:47  */
  assign n15136 = n15093[57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:89:36  */
  assign n15137 = n15135 | n15136;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:72:3  */
  assign n15139 = shifter[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:89:9  */
  assign n15140 = n15137 ? 1'b0 : n15139;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:87:9  */
  assign n15141 = valid_cmd ? 1'b1 : n15140;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:96:24  */
  assign n15142 = shifter[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:97:61  */
  assign n15143 = shifter[8:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:97:66  */
  assign n15145 = n15143 - 5'b00001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:98:31  */
  assign n15146 = n15093[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:98:35  */
  assign n15147 = ~n15146;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:99:41  */
  assign n15148 = shifter[39:9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:99:72  */
  assign n15150 = {n15148, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:101:42  */
  assign n15151 = shifter[40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:101:83  */
  assign n15152 = n15093[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:101:62  */
  assign n15153 = n15151 & n15152;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:101:103  */
  assign n15154 = shifter[40:10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:101:89  */
  assign n15155 = {n15153, n15154};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:98:11  */
  assign n15156 = n15147 ? n15150 : n15155;
  assign n15157 = {n15156, n15145};
  assign n15158 = shifter[40:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:96:9  */
  assign n15159 = n15142 ? n15157 : n15158;
  assign n15160 = {rs1_i, shamt_i};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:93:9  */
  assign n15161 = valid_cmd ? n15160 : n15159;
  assign n15162 = {n15161, n15133};
  assign n15167 = {32'b00000000000000000000000000000000, 5'b00000, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15178 = shifter[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15180 = 1'b0 | n15178;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15182 = shifter[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15183 = n15180 | n15182;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15184 = shifter[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15185 = n15183 | n15184;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15186 = shifter[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15187 = n15185 | n15186;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15188 = shifter[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15189 = n15187 | n15188;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15197 = shifter[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15199 = 1'b0 | n15197;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15201 = shifter[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15202 = n15199 | n15201;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15203 = shifter[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15204 = n15202 | n15203;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n15205 = shifter[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n15206 = n15204 | n15205;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:109:21  */
  assign n15207 = ~n15206;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:110:29  */
  assign n15208 = shifter[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:110:46  */
  assign n15209 = shifter[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:110:34  */
  assign n15210 = n15208 & n15209;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:111:29  */
  assign n15211 = shifter[40:9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:111:48  */
  assign n15212 = shifter[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:111:34  */
  assign n15213 = n15212 ? n15211 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:84:7  */
  always @(posedge clk_i or posedge n15125)
    if (n15125)
      n15215 <= n15167;
    else
      n15215 <= n15162;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:84:7  */
  always @(posedge clk_i or posedge n15125)
    if (n15125)
      n15216 <= 1'b0;
    else
      n15216 <= n15141;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_cp_shifter.vhd:79:7  */
  assign n15217 = {n15215, n15207, n15189, n15216};
endmodule

module neorv32_cpu_decompressor
  (input  [15:0] instr_i,
   output [31:0] instr_o);
  wire illegal;
  wire [31:0] decoded;
  wire n14539;
  wire [3:0] n14545;
  wire [3:0] n14546;
  wire [1:0] n14547;
  wire [9:0] n14548;
  wire n14550;
  wire [10:0] n14551;
  wire [1:0] n14552;
  wire [12:0] n14553;
  wire n14554;
  wire [13:0] n14555;
  wire n14556;
  wire [14:0] n14557;
  wire n14558;
  wire [15:0] n14559;
  wire n14560;
  wire [16:0] n14561;
  wire [2:0] n14562;
  wire [19:0] n14563;
  wire [20:0] n14565;
  wire n14567;
  wire [3:0] n14573;
  wire [4:0] n14574;
  wire [1:0] n14576;
  wire [6:0] n14577;
  wire n14578;
  wire [7:0] n14579;
  wire [1:0] n14580;
  wire [9:0] n14581;
  wire [1:0] n14582;
  wire [11:0] n14583;
  wire [12:0] n14585;
  wire [1:0] n14586;
  wire [2:0] n14587;
  wire [2:0] n14590;
  wire [4:0] n14592;
  wire [3:0] n14594;
  wire [5:0] n14596;
  wire [1:0] n14597;
  wire [7:0] n14598;
  wire n14599;
  wire [8:0] n14600;
  wire n14601;
  wire [9:0] n14602;
  wire [11:0] n14604;
  wire [7:0] n14605;
  wire n14607;
  wire n14610;
  wire n14612;
  wire n14614;
  wire [5:0] n14616;
  wire [2:0] n14617;
  wire [8:0] n14618;
  wire n14619;
  wire [9:0] n14620;
  wire [11:0] n14622;
  wire [2:0] n14624;
  wire [4:0] n14626;
  wire [2:0] n14627;
  wire [4:0] n14629;
  wire n14631;
  wire n14633;
  wire [5:0] n14635;
  wire n14636;
  wire [6:0] n14637;
  wire [1:0] n14638;
  wire n14639;
  wire [2:0] n14640;
  wire [4:0] n14642;
  wire [2:0] n14644;
  wire [4:0] n14646;
  wire [2:0] n14647;
  wire [4:0] n14649;
  wire n14651;
  wire [2:0] n14652;
  reg n14655;
  reg [6:0] n14657;
  reg [4:0] n14659;
  reg [2:0] n14661;
  reg [4:0] n14663;
  wire [4:0] n14664;
  wire [4:0] n14665;
  reg [4:0] n14667;
  wire [6:0] n14668;
  wire [6:0] n14669;
  reg [6:0] n14671;
  wire n14673;
  wire [2:0] n14674;
  wire n14675;
  wire [4:0] n14678;
  wire n14680;
  wire [9:0] n14681;
  wire [10:0] n14682;
  wire n14683;
  wire [11:0] n14684;
  wire [7:0] n14685;
  wire [19:0] n14686;
  wire n14688;
  wire n14690;
  wire n14691;
  wire n14692;
  wire n14693;
  wire [2:0] n14696;
  wire [2:0] n14698;
  wire [4:0] n14700;
  wire n14702;
  wire [5:0] n14703;
  wire [6:0] n14704;
  wire [3:0] n14705;
  wire n14706;
  wire [4:0] n14707;
  wire n14709;
  wire n14711;
  wire n14712;
  wire [4:0] n14714;
  wire n14716;
  wire [3:0] n14722;
  wire [1:0] n14723;
  wire [5:0] n14724;
  wire n14726;
  wire [6:0] n14727;
  wire [4:0] n14728;
  wire [11:0] n14729;
  wire n14731;
  wire [4:0] n14732;
  wire n14734;
  wire n14739;
  wire [2:0] n14745;
  wire [1:0] n14747;
  wire [4:0] n14748;
  wire n14749;
  wire [5:0] n14750;
  wire n14751;
  wire [6:0] n14752;
  wire n14753;
  wire [7:0] n14754;
  wire [11:0] n14756;
  wire [4:0] n14758;
  wire n14760;
  wire [3:0] n14766;
  wire [3:0] n14767;
  wire [3:0] n14768;
  wire [2:0] n14769;
  wire [14:0] n14770;
  wire [4:0] n14772;
  wire [19:0] n14773;
  wire [31:0] n14774;
  wire [31:0] n14775;
  wire [31:0] n14776;
  wire [4:0] n14777;
  wire n14779;
  wire n14780;
  wire n14781;
  wire n14782;
  wire n14785;
  wire n14787;
  wire [4:0] n14788;
  wire [4:0] n14789;
  wire n14791;
  wire [3:0] n14797;
  wire [2:0] n14798;
  wire [6:0] n14799;
  wire [4:0] n14801;
  wire [11:0] n14802;
  wire n14804;
  wire [2:0] n14805;
  wire [4:0] n14807;
  wire [2:0] n14808;
  wire [4:0] n14810;
  wire [2:0] n14811;
  wire [4:0] n14813;
  wire [1:0] n14814;
  wire n14815;
  wire n14816;
  wire [6:0] n14819;
  wire [4:0] n14821;
  wire n14822;
  wire n14825;
  wire n14827;
  wire n14829;
  wire n14830;
  wire n14833;
  wire [3:0] n14839;
  wire [2:0] n14840;
  wire [6:0] n14841;
  wire [4:0] n14843;
  wire [11:0] n14844;
  wire n14846;
  wire [1:0] n14848;
  wire n14851;
  wire n14855;
  wire n14859;
  wire [2:0] n14861;
  reg [2:0] n14862;
  reg [6:0] n14863;
  wire n14864;
  wire n14867;
  wire [1:0] n14868;
  reg n14870;
  reg [6:0] n14871;
  reg [2:0] n14872;
  wire [4:0] n14873;
  reg [4:0] n14874;
  wire [6:0] n14875;
  reg [6:0] n14876;
  wire [4:0] n14877;
  reg n14879;
  wire [6:0] n14880;
  reg [6:0] n14881;
  wire [4:0] n14882;
  reg [4:0] n14883;
  wire [2:0] n14884;
  wire [2:0] n14885;
  reg [2:0] n14886;
  wire [4:0] n14887;
  wire [4:0] n14888;
  reg [4:0] n14889;
  wire [4:0] n14890;
  wire [4:0] n14891;
  wire [4:0] n14892;
  wire [4:0] n14893;
  reg [4:0] n14894;
  wire [6:0] n14895;
  wire [6:0] n14896;
  wire [6:0] n14897;
  wire [6:0] n14898;
  reg [6:0] n14899;
  wire n14901;
  wire [2:0] n14902;
  wire [4:0] n14903;
  wire [4:0] n14904;
  wire [4:0] n14907;
  wire n14908;
  wire n14911;
  wire n14913;
  wire [1:0] n14914;
  wire [5:0] n14916;
  wire n14917;
  wire [6:0] n14918;
  wire [2:0] n14919;
  wire [9:0] n14920;
  wire [11:0] n14922;
  wire [4:0] n14924;
  wire n14925;
  wire [4:0] n14926;
  wire n14928;
  wire n14929;
  wire n14932;
  wire n14934;
  wire n14936;
  wire n14937;
  wire [1:0] n14938;
  wire [5:0] n14940;
  wire n14941;
  wire [6:0] n14942;
  wire [2:0] n14943;
  wire [4:0] n14945;
  wire [4:0] n14947;
  wire n14948;
  wire n14951;
  wire n14953;
  wire n14955;
  wire n14956;
  wire n14957;
  wire n14958;
  wire [4:0] n14959;
  wire n14961;
  wire [4:0] n14963;
  wire [4:0] n14965;
  wire n14967;
  wire [4:0] n14968;
  wire n14970;
  wire n14971;
  wire n14974;
  wire [4:0] n14976;
  wire [4:0] n14978;
  wire [4:0] n14979;
  wire n14981;
  wire n14984;
  wire n14985;
  wire [24:0] n14986;
  wire [11:0] n14987;
  wire [11:0] n14988;
  wire [11:0] n14989;
  wire [2:0] n14990;
  wire [2:0] n14992;
  wire [4:0] n14993;
  wire [4:0] n14994;
  wire [4:0] n14995;
  wire [4:0] n14997;
  wire [4:0] n14998;
  wire n15000;
  wire [4:0] n15001;
  wire n15003;
  wire [4:0] n15006;
  wire [11:0] n15008;
  wire [6:0] n15009;
  wire [6:0] n15010;
  wire [4:0] n15011;
  wire [4:0] n15013;
  wire [4:0] n15015;
  wire [11:0] n15017;
  wire [4:0] n15019;
  wire [4:0] n15020;
  wire [4:0] n15021;
  wire [24:0] n15022;
  wire [11:0] n15023;
  wire [16:0] n15024;
  wire [11:0] n15025;
  wire [11:0] n15026;
  wire [2:0] n15027;
  wire [2:0] n15029;
  wire [9:0] n15030;
  wire [9:0] n15031;
  wire [9:0] n15032;
  wire [6:0] n15033;
  wire [6:0] n15035;
  wire n15037;
  wire [31:0] n15038;
  wire [24:0] n15039;
  wire [24:0] n15040;
  wire [24:0] n15041;
  wire [6:0] n15042;
  wire [6:0] n15044;
  wire n15046;
  wire [3:0] n15047;
  reg n15049;
  wire [6:0] n15050;
  reg [6:0] n15052;
  wire [4:0] n15053;
  reg [4:0] n15055;
  wire [2:0] n15056;
  reg [2:0] n15058;
  wire [4:0] n15059;
  reg [4:0] n15061;
  wire [4:0] n15062;
  wire [4:0] n15063;
  reg [4:0] n15065;
  wire [6:0] n15066;
  reg [6:0] n15068;
  wire [1:0] n15069;
  reg n15070;
  reg [6:0] n15072;
  reg [4:0] n15073;
  reg [2:0] n15074;
  reg [4:0] n15075;
  reg [4:0] n15076;
  reg [6:0] n15077;
  wire [29:0] n15085;
  wire n15086;
  wire n15087;
  wire n15088;
  wire n15090;
  wire [31:0] n15091;
  wire [31:0] n15092;
  assign instr_o = n15092; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:45:10  */
  assign illegal = n15070; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:46:10  */
  assign decoded = n15091; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:35  */
  assign n14539 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:175:9  */
  assign n14545 = {n14539, n14539, n14539, n14539};
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:177:22  */
  assign n14546 = {n14539, n14539, n14539, n14539};
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:173:7  */
  assign n14547 = {n14539, n14539};
  assign n14548 = {n14545, n14546, n14547};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:53  */
  assign n14550 = instr_i[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:44  */
  assign n14551 = {n14548, n14550};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:66  */
  assign n14552 = instr_i[10:9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:57  */
  assign n14553 = {n14551, n14552};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:89  */
  assign n14554 = instr_i[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:80  */
  assign n14555 = {n14553, n14554};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:102  */
  assign n14556 = instr_i[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:93  */
  assign n14557 = {n14555, n14556};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:115  */
  assign n14558 = instr_i[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:106  */
  assign n14559 = {n14557, n14558};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:128  */
  assign n14560 = instr_i[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:119  */
  assign n14561 = {n14559, n14560};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:142  */
  assign n14562 = instr_i[5:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:133  */
  assign n14563 = {n14561, n14562};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:57:155  */
  assign n14565 = {n14563, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:35  */
  assign n14567 = instr_i[12]; // extract
  assign n14573 = {n14567, n14567, n14567, n14567};
  assign n14574 = {n14573, n14567};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:52  */
  assign n14576 = instr_i[6:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:43  */
  assign n14577 = {n14574, n14576};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:74  */
  assign n14578 = instr_i[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:65  */
  assign n14579 = {n14577, n14578};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:87  */
  assign n14580 = instr_i[11:10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:78  */
  assign n14581 = {n14579, n14580};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:111  */
  assign n14582 = instr_i[4:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:102  */
  assign n14583 = {n14581, n14582};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:58:124  */
  assign n14585 = {n14583, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:65:17  */
  assign n14586 = instr_i[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:68:21  */
  assign n14587 = instr_i[15:13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:74:84  */
  assign n14590 = instr_i[4:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:74:75  */
  assign n14592 = {2'b01, n14590};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:84  */
  assign n14594 = instr_i[10:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:75  */
  assign n14596 = {2'b00, n14594};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:107  */
  assign n14597 = instr_i[12:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:98  */
  assign n14598 = {n14596, n14597};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:131  */
  assign n14599 = instr_i[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:122  */
  assign n14600 = {n14598, n14599};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:144  */
  assign n14601 = instr_i[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:135  */
  assign n14602 = {n14600, n14601};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:76:148  */
  assign n14604 = {n14602, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:77:24  */
  assign n14605 = instr_i[12:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:77:38  */
  assign n14607 = n14605 == 8'b00000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:77:13  */
  assign n14610 = n14607 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:70:11  */
  assign n14612 = n14587 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:84:87  */
  assign n14614 = instr_i[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:84:78  */
  assign n14616 = {5'b00000, n14614};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:84:100  */
  assign n14617 = instr_i[12:10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:84:91  */
  assign n14618 = {n14616, n14617};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:84:124  */
  assign n14619 = instr_i[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:84:115  */
  assign n14620 = {n14618, n14619};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:84:128  */
  assign n14622 = {n14620, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:86:84  */
  assign n14624 = instr_i[9:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:86:75  */
  assign n14626 = {2'b01, n14624};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:87:84  */
  assign n14627 = instr_i[4:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:87:75  */
  assign n14629 = {2'b01, n14627};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:81:11  */
  assign n14631 = n14587 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:92:87  */
  assign n14633 = instr_i[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:92:78  */
  assign n14635 = {5'b00000, n14633};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:92:100  */
  assign n14636 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:92:91  */
  assign n14637 = {n14635, n14636};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:93:77  */
  assign n14638 = instr_i[11:10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:93:101  */
  assign n14639 = instr_i[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:93:92  */
  assign n14640 = {n14638, n14639};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:93:105  */
  assign n14642 = {n14640, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:95:84  */
  assign n14644 = instr_i[9:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:95:75  */
  assign n14646 = {2'b01, n14644};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:96:84  */
  assign n14647 = instr_i[4:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:96:75  */
  assign n14649 = {2'b01, n14647};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:89:11  */
  assign n14651 = n14587 == 3'b110;
  assign n14652 = {n14651, n14631, n14612};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:68:9  */
  always @*
    case (n14652)
      3'b100: n14655 = 1'b0;
      3'b010: n14655 = 1'b0;
      3'b001: n14655 = n14610;
      default: n14655 = 1'b1;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:68:9  */
  always @*
    case (n14652)
      3'b100: n14657 = 7'b0100011;
      3'b010: n14657 = 7'b0000011;
      3'b001: n14657 = 7'b0010011;
      default: n14657 = 7'b0000011;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:68:9  */
  always @*
    case (n14652)
      3'b100: n14659 = n14642;
      3'b010: n14659 = n14629;
      3'b001: n14659 = n14592;
      default: n14659 = 5'b00000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:68:9  */
  always @*
    case (n14652)
      3'b100: n14661 = 3'b010;
      3'b010: n14661 = 3'b010;
      3'b001: n14661 = 3'b000;
      default: n14661 = 3'b000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:68:9  */
  always @*
    case (n14652)
      3'b100: n14663 = n14646;
      3'b010: n14663 = n14626;
      3'b001: n14663 = 5'b00010;
      default: n14663 = 5'b00000;
    endcase
  assign n14664 = n14604[4:0]; // extract
  assign n14665 = n14622[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:68:9  */
  always @*
    case (n14652)
      3'b100: n14667 = n14649;
      3'b010: n14667 = n14665;
      3'b001: n14667 = n14664;
      default: n14667 = 5'b00000;
    endcase
  assign n14668 = n14604[11:5]; // extract
  assign n14669 = n14622[11:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:68:9  */
  always @*
    case (n14652)
      3'b100: n14671 = n14637;
      3'b010: n14671 = n14669;
      3'b001: n14671 = n14668;
      default: n14671 = 7'b0000000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:67:7  */
  assign n14673 = n14586 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:21  */
  assign n14674 = instr_i[15:13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:110:24  */
  assign n14675 = instr_i[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:110:13  */
  assign n14678 = n14675 ? 5'b00000 : 5'b00001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:116:77  */
  assign n14680 = n14565[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:116:91  */
  assign n14681 = n14565[10:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:116:82  */
  assign n14682 = {n14680, n14681};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:116:114  */
  assign n14683 = n14565[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:116:105  */
  assign n14684 = {n14682, n14683};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:116:128  */
  assign n14685 = n14565[19:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:116:119  */
  assign n14686 = {n14684, n14685};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:108:11  */
  assign n14688 = n14674 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:108:22  */
  assign n14690 = n14674 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:108:22  */
  assign n14691 = n14688 | n14690;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:120:24  */
  assign n14692 = instr_i[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:120:42  */
  assign n14693 = ~n14692;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:120:13  */
  assign n14696 = n14693 ? 3'b000 : 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:126:84  */
  assign n14698 = instr_i[9:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:126:75  */
  assign n14700 = {2'b01, n14698};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:128:77  */
  assign n14702 = n14585[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:128:91  */
  assign n14703 = n14585[10:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:128:82  */
  assign n14704 = {n14702, n14703};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:129:77  */
  assign n14705 = n14585[4:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:129:99  */
  assign n14706 = n14585[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:129:90  */
  assign n14707 = {n14705, n14706};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:11  */
  assign n14709 = n14674 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:22  */
  assign n14711 = n14674 == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:118:22  */
  assign n14712 = n14709 | n14711;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:136:77  */
  assign n14714 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:137:89  */
  assign n14716 = instr_i[12]; // extract
  assign n14722 = {n14716, n14716, n14716, n14716};
  assign n14723 = {n14716, n14716};
  assign n14724 = {n14722, n14723};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:137:106  */
  assign n14726 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:137:97  */
  assign n14727 = {n14724, n14726};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:137:120  */
  assign n14728 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:137:111  */
  assign n14729 = {n14727, n14728};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:131:11  */
  assign n14731 = n14674 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:141:24  */
  assign n14732 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:141:61  */
  assign n14734 = n14732 == 5'b00010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:91  */
  assign n14739 = instr_i[12]; // extract
  assign n14745 = {n14739, n14739, n14739};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:108  */
  assign n14747 = instr_i[4:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:99  */
  assign n14748 = {n14745, n14747};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:130  */
  assign n14749 = instr_i[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:121  */
  assign n14750 = {n14748, n14749};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:143  */
  assign n14751 = instr_i[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:134  */
  assign n14752 = {n14750, n14751};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:156  */
  assign n14753 = instr_i[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:147  */
  assign n14754 = {n14752, n14753};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:147:160  */
  assign n14756 = {n14754, 4'b0000};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:150:79  */
  assign n14758 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:151:91  */
  assign n14760 = instr_i[12]; // extract
  assign n14766 = {n14760, n14760, n14760, n14760};
  assign n14767 = {n14760, n14760, n14760, n14760};
  assign n14768 = {n14760, n14760, n14760, n14760};
  assign n14769 = {n14760, n14760, n14760};
  assign n14770 = {n14766, n14767, n14768, n14769};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:151:109  */
  assign n14772 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:151:100  */
  assign n14773 = {n14770, n14772};
  assign n14774 = {n14773, n14758, 7'b0110111};
  assign n14775 = {n14756, 5'b00010, 3'b000, 5'b00010, 7'b0010011};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:141:13  */
  assign n14776 = n14734 ? n14775 : n14774;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:153:24  */
  assign n14777 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:153:37  */
  assign n14779 = n14777 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:153:60  */
  assign n14780 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:153:65  */
  assign n14781 = ~n14780;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:153:48  */
  assign n14782 = n14781 & n14779;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:153:13  */
  assign n14785 = n14782 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:139:11  */
  assign n14787 = n14674 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:161:77  */
  assign n14788 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:162:77  */
  assign n14789 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:163:89  */
  assign n14791 = instr_i[12]; // extract
  assign n14797 = {n14791, n14791, n14791, n14791};
  assign n14798 = {n14791, n14791, n14791};
  assign n14799 = {n14797, n14798};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:163:106  */
  assign n14801 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:163:97  */
  assign n14802 = {n14799, n14801};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:157:11  */
  assign n14804 = n14674 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:167:78  */
  assign n14805 = instr_i[9:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:167:69  */
  assign n14807 = {2'b01, n14805};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:168:78  */
  assign n14808 = instr_i[9:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:168:69  */
  assign n14810 = {2'b01, n14808};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:169:78  */
  assign n14811 = instr_i[4:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:169:69  */
  assign n14813 = {2'b01, n14811};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:170:25  */
  assign n14814 = instr_i[11:10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:172:28  */
  assign n14815 = instr_i[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:172:33  */
  assign n14816 = ~n14815;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:172:17  */
  assign n14819 = n14816 ? 7'b0000000 : 7'b0100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:179:81  */
  assign n14821 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:180:28  */
  assign n14822 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:180:17  */
  assign n14825 = n14822 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:171:15  */
  assign n14827 = n14814 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:171:25  */
  assign n14829 = n14814 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:171:25  */
  assign n14830 = n14827 | n14829;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:186:93  */
  assign n14833 = instr_i[12]; // extract
  assign n14839 = {n14833, n14833, n14833, n14833};
  assign n14840 = {n14833, n14833, n14833};
  assign n14841 = {n14839, n14840};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:186:110  */
  assign n14843 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:186:101  */
  assign n14844 = {n14841, n14843};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:183:15  */
  assign n14846 = n14814 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:189:29  */
  assign n14848 = instr_i[6:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:190:19  */
  assign n14851 = n14848 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:193:19  */
  assign n14855 = n14848 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:196:19  */
  assign n14859 = n14848 == 2'b10;
  assign n14861 = {n14859, n14855, n14851};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:189:17  */
  always @*
    case (n14861)
      3'b100: n14862 = 3'b110;
      3'b010: n14862 = 3'b100;
      3'b001: n14862 = 3'b000;
      default: n14862 = 3'b111;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:189:17  */
  always @*
    case (n14861)
      3'b100: n14863 = 7'b0000000;
      3'b010: n14863 = 7'b0000000;
      3'b001: n14863 = 7'b0100000;
      default: n14863 = 7'b0000000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:203:28  */
  assign n14864 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:203:17  */
  assign n14867 = n14864 ? 1'b1 : 1'b0;
  assign n14868 = {n14846, n14830};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:170:13  */
  always @*
    case (n14868)
      2'b10: n14870 = 1'b0;
      2'b01: n14870 = n14825;
      default: n14870 = n14867;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:170:13  */
  always @*
    case (n14868)
      2'b10: n14871 = 7'b0010011;
      2'b01: n14871 = 7'b0010011;
      default: n14871 = 7'b0110011;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:170:13  */
  always @*
    case (n14868)
      2'b10: n14872 = 3'b111;
      2'b01: n14872 = 3'b101;
      default: n14872 = n14862;
    endcase
  assign n14873 = n14844[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:170:13  */
  always @*
    case (n14868)
      2'b10: n14874 = n14873;
      2'b01: n14874 = n14821;
      default: n14874 = n14813;
    endcase
  assign n14875 = n14844[11:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:170:13  */
  always @*
    case (n14868)
      2'b10: n14876 = n14875;
      2'b01: n14876 = n14819;
      default: n14876 = n14863;
    endcase
  assign n14877 = {n14804, n14787, n14731, n14712, n14691};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:9  */
  always @*
    case (n14877)
      5'b10000: n14879 = 1'b0;
      5'b01000: n14879 = n14785;
      5'b00100: n14879 = 1'b0;
      5'b00010: n14879 = 1'b0;
      5'b00001: n14879 = 1'b0;
      default: n14879 = n14870;
    endcase
  assign n14880 = n14776[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:9  */
  always @*
    case (n14877)
      5'b10000: n14881 = 7'b0010011;
      5'b01000: n14881 = n14880;
      5'b00100: n14881 = 7'b0010011;
      5'b00010: n14881 = 7'b1100011;
      5'b00001: n14881 = 7'b1101111;
      default: n14881 = n14871;
    endcase
  assign n14882 = n14776[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:9  */
  always @*
    case (n14877)
      5'b10000: n14883 = n14789;
      5'b01000: n14883 = n14882;
      5'b00100: n14883 = n14714;
      5'b00010: n14883 = n14707;
      5'b00001: n14883 = n14678;
      default: n14883 = n14807;
    endcase
  assign n14884 = n14686[2:0]; // extract
  assign n14885 = n14776[14:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:9  */
  always @*
    case (n14877)
      5'b10000: n14886 = 3'b000;
      5'b01000: n14886 = n14885;
      5'b00100: n14886 = 3'b000;
      5'b00010: n14886 = n14696;
      5'b00001: n14886 = n14884;
      default: n14886 = n14872;
    endcase
  assign n14887 = n14686[7:3]; // extract
  assign n14888 = n14776[19:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:9  */
  always @*
    case (n14877)
      5'b10000: n14889 = n14788;
      5'b01000: n14889 = n14888;
      5'b00100: n14889 = 5'b00000;
      5'b00010: n14889 = n14700;
      5'b00001: n14889 = n14887;
      default: n14889 = n14810;
    endcase
  assign n14890 = n14686[12:8]; // extract
  assign n14891 = n14729[4:0]; // extract
  assign n14892 = n14776[24:20]; // extract
  assign n14893 = n14802[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:9  */
  always @*
    case (n14877)
      5'b10000: n14894 = n14893;
      5'b01000: n14894 = n14892;
      5'b00100: n14894 = n14891;
      5'b00010: n14894 = 5'b00000;
      5'b00001: n14894 = n14890;
      default: n14894 = n14874;
    endcase
  assign n14895 = n14686[19:13]; // extract
  assign n14896 = n14729[11:5]; // extract
  assign n14897 = n14776[31:25]; // extract
  assign n14898 = n14802[11:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:106:9  */
  always @*
    case (n14877)
      5'b10000: n14899 = n14898;
      5'b01000: n14899 = n14897;
      5'b00100: n14899 = n14896;
      5'b00010: n14899 = n14704;
      5'b00001: n14899 = n14895;
      default: n14899 = n14876;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:104:7  */
  assign n14901 = n14586 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:211:21  */
  assign n14902 = instr_i[15:13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:216:77  */
  assign n14903 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:217:77  */
  assign n14904 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:220:77  */
  assign n14907 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:221:24  */
  assign n14908 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:221:13  */
  assign n14911 = n14908 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:213:11  */
  assign n14913 = n14902 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:86  */
  assign n14914 = instr_i[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:77  */
  assign n14916 = {4'b0000, n14914};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:108  */
  assign n14917 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:99  */
  assign n14918 = {n14916, n14917};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:122  */
  assign n14919 = instr_i[6:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:113  */
  assign n14920 = {n14918, n14919};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:228:135  */
  assign n14922 = {n14920, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:231:77  */
  assign n14924 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:232:24  */
  assign n14925 = instr_i[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:233:24  */
  assign n14926 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:233:61  */
  assign n14928 = n14926 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:232:49  */
  assign n14929 = n14925 | n14928;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:232:13  */
  assign n14932 = n14929 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:225:11  */
  assign n14934 = n14902 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:225:22  */
  assign n14936 = n14902 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:225:22  */
  assign n14937 = n14934 | n14936;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:240:86  */
  assign n14938 = instr_i[8:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:240:77  */
  assign n14940 = {4'b0000, n14938};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:240:108  */
  assign n14941 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:240:99  */
  assign n14942 = {n14940, n14941};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:241:77  */
  assign n14943 = instr_i[11:9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:241:91  */
  assign n14945 = {n14943, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:244:77  */
  assign n14947 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:245:24  */
  assign n14948 = instr_i[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:245:13  */
  assign n14951 = n14948 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:237:11  */
  assign n14953 = n14902 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:237:22  */
  assign n14955 = n14902 == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:237:22  */
  assign n14956 = n14953 | n14955;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:251:24  */
  assign n14957 = instr_i[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:251:29  */
  assign n14958 = ~n14957;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:252:26  */
  assign n14959 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:252:39  */
  assign n14961 = n14959 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:254:81  */
  assign n14963 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:28  */
  assign n14965 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:67  */
  assign n14967 = n14965 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:257:28  */
  assign n14968 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:257:67  */
  assign n14970 = n14968 != 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:78  */
  assign n14971 = n14967 | n14970;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:256:17  */
  assign n14974 = n14971 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:263:81  */
  assign n14976 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:265:81  */
  assign n14978 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:28  */
  assign n14979 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:67  */
  assign n14981 = n14979 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:266:17  */
  assign n14984 = n14981 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:252:15  */
  assign n14985 = n14961 ? n14974 : n14984;
  assign n14986 = {n14978, 5'b00000, 3'b000, n14976, 7'b0110011};
  assign n14987 = {5'b00000, 7'b1100111};
  assign n14988 = n14986[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:252:15  */
  assign n14989 = n14961 ? n14987 : n14988;
  assign n14990 = n14986[14:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:252:15  */
  assign n14992 = n14961 ? 3'b000 : n14990;
  assign n14993 = n14986[19:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:252:15  */
  assign n14994 = n14961 ? n14963 : n14993;
  assign n14995 = n14986[24:20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:252:15  */
  assign n14997 = n14961 ? 5'b00000 : n14995;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:271:26  */
  assign n14998 = instr_i[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:271:39  */
  assign n15000 = n14998 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:272:28  */
  assign n15001 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:272:42  */
  assign n15003 = n15001 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:277:83  */
  assign n15006 = instr_i[11:7]; // extract
  assign n15008 = {5'b00001, 7'b1100111};
  assign n15009 = n15008[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:272:17  */
  assign n15010 = n15003 ? 7'b1110011 : n15009;
  assign n15011 = n15008[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:272:17  */
  assign n15013 = n15003 ? 5'b00000 : n15011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:272:17  */
  assign n15015 = n15003 ? 5'b00000 : n15006;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:272:17  */
  assign n15017 = n15003 ? 12'b000000000001 : 12'b000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:283:81  */
  assign n15019 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:284:81  */
  assign n15020 = instr_i[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:285:81  */
  assign n15021 = instr_i[6:2]; // extract
  assign n15022 = {n15021, n15020, 3'b000, n15019, 7'b0110011};
  assign n15023 = {n15013, n15010};
  assign n15024 = {n15017, n15015};
  assign n15025 = n15022[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:271:15  */
  assign n15026 = n15000 ? n15023 : n15025;
  assign n15027 = n15022[14:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:271:15  */
  assign n15029 = n15000 ? 3'b000 : n15027;
  assign n15030 = n15022[24:15]; // extract
  assign n15031 = n15024[9:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:271:15  */
  assign n15032 = n15000 ? n15031 : n15030;
  assign n15033 = n15024[16:10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:271:15  */
  assign n15035 = n15000 ? n15033 : 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:251:13  */
  assign n15037 = n14958 ? n14985 : 1'b0;
  assign n15038 = {n15035, n15032, n15029, n15026};
  assign n15039 = {n14997, n14994, n14992, n14989};
  assign n15040 = n15038[24:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:251:13  */
  assign n15041 = n14958 ? n15039 : n15040;
  assign n15042 = n15038[31:25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:251:13  */
  assign n15044 = n14958 ? 7'b0000000 : n15042;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:249:11  */
  assign n15046 = n14902 == 3'b100;
  assign n15047 = {n15046, n14956, n14937, n14913};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:211:9  */
  always @*
    case (n15047)
      4'b1000: n15049 = n15037;
      4'b0100: n15049 = n14951;
      4'b0010: n15049 = n14932;
      4'b0001: n15049 = n14911;
      default: n15049 = 1'b1;
    endcase
  assign n15050 = n15041[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:211:9  */
  always @*
    case (n15047)
      4'b1000: n15052 = n15050;
      4'b0100: n15052 = 7'b0100011;
      4'b0010: n15052 = 7'b0000011;
      4'b0001: n15052 = 7'b0010011;
      default: n15052 = 7'b0000011;
    endcase
  assign n15053 = n15041[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:211:9  */
  always @*
    case (n15047)
      4'b1000: n15055 = n15053;
      4'b0100: n15055 = n14945;
      4'b0010: n15055 = n14924;
      4'b0001: n15055 = n14904;
      default: n15055 = 5'b00000;
    endcase
  assign n15056 = n15041[14:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:211:9  */
  always @*
    case (n15047)
      4'b1000: n15058 = n15056;
      4'b0100: n15058 = 3'b010;
      4'b0010: n15058 = 3'b010;
      4'b0001: n15058 = 3'b001;
      default: n15058 = 3'b000;
    endcase
  assign n15059 = n15041[19:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:211:9  */
  always @*
    case (n15047)
      4'b1000: n15061 = n15059;
      4'b0100: n15061 = 5'b00010;
      4'b0010: n15061 = 5'b00010;
      4'b0001: n15061 = n14903;
      default: n15061 = 5'b00000;
    endcase
  assign n15062 = n14922[4:0]; // extract
  assign n15063 = n15041[24:20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:211:9  */
  always @*
    case (n15047)
      4'b1000: n15065 = n15063;
      4'b0100: n15065 = n14947;
      4'b0010: n15065 = n15062;
      4'b0001: n15065 = n14907;
      default: n15065 = 5'b00000;
    endcase
  assign n15066 = n14922[11:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:211:9  */
  always @*
    case (n15047)
      4'b1000: n15068 = n15044;
      4'b0100: n15068 = n14942;
      4'b0010: n15068 = n15066;
      4'b0001: n15068 = 7'b0000000;
      default: n15068 = 7'b0000000;
    endcase
  assign n15069 = {n14901, n14673};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:65:5  */
  always @*
    case (n15069)
      2'b10: n15070 = n14879;
      2'b01: n15070 = n14655;
      default: n15070 = n15049;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:65:5  */
  always @*
    case (n15069)
      2'b10: n15072 = n14881;
      2'b01: n15072 = n14657;
      default: n15072 = n15052;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:65:5  */
  always @*
    case (n15069)
      2'b10: n15073 = n14883;
      2'b01: n15073 = n14659;
      default: n15073 = n15055;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:65:5  */
  always @*
    case (n15069)
      2'b10: n15074 = n14886;
      2'b01: n15074 = n14661;
      default: n15074 = n15058;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:65:5  */
  always @*
    case (n15069)
      2'b10: n15075 = n14889;
      2'b01: n15075 = n14663;
      default: n15075 = n15061;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:65:5  */
  always @*
    case (n15069)
      2'b10: n15076 = n14894;
      2'b01: n15076 = n14667;
      default: n15076 = n15065;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:65:5  */
  always @*
    case (n15069)
      2'b10: n15077 = n14899;
      2'b01: n15077 = n14671;
      default: n15077 = n15068;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:299:34  */
  assign n15085 = decoded[31:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:300:24  */
  assign n15086 = decoded[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:300:42  */
  assign n15087 = ~illegal;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:300:28  */
  assign n15088 = n15087 ? n15086 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_decompressor.vhd:301:24  */
  assign n15090 = decoded[0]; // extract
  assign n15091 = {n15077, n15076, n15075, n15074, n15073, n15072};
  assign n15092 = {n15085, n15088, n15090};
endmodule

module neorv32_fifo_2_17_29e2dcfbb16f63bb0254df7585a15bb6fb5e927d
  (input  clk_i,
   input  rstn_i,
   input  clear_i,
   input  [16:0] wdata_i,
   input  we_i,
   input  re_i,
   output half_o,
   output free_o,
   output [16:0] rdata_o,
   output avail_o);
  wire we;
  wire re;
  wire match;
  wire empty;
  wire full;
  wire half;
  wire free;
  wire avail;
  wire [1:0] w_pnt;
  wire [1:0] w_nxt;
  wire [1:0] r_pnt;
  wire [1:0] r_nxt;
  wire [1:0] r_pnt_ff;
  wire [1:0] diff;
  wire n14455;
  wire n14456;
  wire n14458;
  wire n14459;
  wire n14461;
  wire [1:0] n14471;
  wire [1:0] n14473;
  wire [1:0] n14474;
  wire [1:0] n14476;
  wire [1:0] n14478;
  wire [1:0] n14479;
  wire n14481;
  wire n14482;
  wire n14483;
  wire n14484;
  wire n14487;
  wire n14488;
  wire n14489;
  wire n14490;
  wire n14491;
  wire n14494;
  wire n14495;
  wire n14496;
  wire n14497;
  wire n14498;
  wire [1:0] n14500;
  wire n14501;
  wire n14502;
  wire n14503;
  wire n14504;
  wire n14507;
  wire n14520;
  reg [1:0] n14529;
  reg [1:0] n14530;
  reg [1:0] n14531;
  wire [16:0] n14532; // mem_rd
  assign half_o = half; //(module output)
  assign free_o = free; //(module output)
  assign rdata_o = n14532; //(module output)
  assign avail_o = avail; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:10  */
  assign we = n14458; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:14  */
  assign re = n14455; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:18  */
  assign match = n14484; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:25  */
  assign empty = n14498; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:32  */
  assign full = n14491; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:38  */
  assign half = n14502; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:44  */
  assign free = n14503; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:50  */
  assign avail = n14504; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:10  */
  assign w_pnt = n14529; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:17  */
  assign w_nxt = n14471; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:24  */
  assign r_pnt = n14530; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:31  */
  assign r_nxt = n14476; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:38  */
  assign r_pnt_ff = n14531; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:60:10  */
  assign diff = n14500; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:66:14  */
  assign n14455 = 1'b1 ? re_i : n14456;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:66:50  */
  assign n14456 = re_i & avail;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:67:14  */
  assign n14458 = 1'b1 ? we_i : n14459;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:67:50  */
  assign n14459 = we_i & free;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:74:16  */
  assign n14461 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:28  */
  assign n14471 = clear_i ? 2'b00 : n14474;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:88  */
  assign n14473 = w_pnt + 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:49  */
  assign n14474 = we ? n14473 : w_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:28  */
  assign n14476 = clear_i ? 2'b00 : n14479;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:88  */
  assign n14478 = r_pnt + 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:49  */
  assign n14479 = re ? n14478 : r_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:94:29  */
  assign n14481 = r_pnt[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:94:60  */
  assign n14482 = w_pnt[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:94:53  */
  assign n14483 = n14481 == n14482;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:94:18  */
  assign n14484 = n14483 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:95:29  */
  assign n14487 = r_pnt[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:95:50  */
  assign n14488 = w_pnt[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:95:42  */
  assign n14489 = n14487 != n14488;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:95:64  */
  assign n14490 = match & n14489;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:95:18  */
  assign n14491 = n14490 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:96:29  */
  assign n14494 = r_pnt[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:96:50  */
  assign n14495 = w_pnt[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:96:43  */
  assign n14496 = n14494 == n14495;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:96:64  */
  assign n14497 = match & n14496;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:96:18  */
  assign n14498 = n14497 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:97:48  */
  assign n14500 = w_pnt - r_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:98:18  */
  assign n14501 = diff[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:98:32  */
  assign n14502 = n14501 | full;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:110:12  */
  assign n14503 = ~full;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:111:12  */
  assign n14504 = ~empty;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:177:47  */
  assign n14507 = w_pnt[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:206:55  */
  assign n14520 = r_pnt_ff[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:77:5  */
  always @(posedge clk_i or posedge n14461)
    if (n14461)
      n14529 <= 2'b00;
    else
      n14529 <= w_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:77:5  */
  always @(posedge clk_i or posedge n14461)
    if (n14461)
      n14530 <= 2'b00;
    else
      n14530 <= r_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:202:9  */
  always @(posedge clk_i)
    n14531 <= r_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:206:27  */
  reg [16:0] fifo_mem[1:0] ; // memory
  assign n14532 = fifo_mem[n14520];
  always @(posedge clk_i)
    if (we)
      fifo_mem[n14507] <= wdata_i;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:206:27  */
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:177:22  */
endmodule

module neorv32_pwm_channel
  (input  clk_i,
   input  rstn_i,
   input  we_i,
   input  re_i,
   input  [31:0] wdata_i,
   input  [7:0] clkgen_i,
   output [31:0] rdata_o,
   output clkgen_en_o,
   output pwm_o);
  wire cfg_en;
  wire [2:0] cfg_prsc;
  wire [9:0] cfg_cdiv;
  wire [7:0] cfg_duty;
  wire [9:0] cnt_cdiv;
  wire cnt_tick;
  wire [7:0] cnt_duty;
  wire n14368;
  wire n14370;
  wire [2:0] n14371;
  wire [9:0] n14372;
  wire [7:0] n14373;
  wire [3:0] n14391;
  wire [13:0] n14393;
  wire [23:0] n14394;
  wire [31:0] n14395;
  wire [31:0] n14396;
  wire n14399;
  wire n14401;
  wire [9:0] n14406;
  wire [9:0] n14408;
  wire [9:0] n14409;
  wire [9:0] n14411;
  wire n14412;
  wire [7:0] n14414;
  wire [7:0] n14415;
  wire [7:0] n14417;
  wire n14418;
  wire n14419;
  wire n14420;
  wire n14423;
  wire n14435;
  wire n14436;
  wire n14438;
  reg n14439;
  wire [2:0] n14440;
  reg [2:0] n14441;
  wire [9:0] n14442;
  reg [9:0] n14443;
  wire [7:0] n14444;
  reg [7:0] n14445;
  reg [9:0] n14446;
  reg [7:0] n14447;
  reg n14448;
  wire n14449;
  assign rdata_o = n14396; //(module output)
  assign clkgen_en_o = cfg_en; //(module output)
  assign pwm_o = n14448; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:159:10  */
  assign cfg_en = n14439; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:160:10  */
  assign cfg_prsc = n14441; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:161:10  */
  assign cfg_cdiv = n14443; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:162:10  */
  assign cfg_duty = n14445; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:165:10  */
  assign cnt_cdiv = n14446; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:166:10  */
  assign cnt_tick = n14436; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:167:10  */
  assign cnt_duty = n14447; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:175:16  */
  assign n14368 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:182:28  */
  assign n14370 = wdata_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:183:28  */
  assign n14371 = wdata_i[30:28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:184:28  */
  assign n14372 = wdata_i[17:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:185:28  */
  assign n14373 = wdata_i[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:191:21  */
  assign n14391 = {cfg_en, cfg_prsc};
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:191:32  */
  assign n14393 = {n14391, 10'b0000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:191:47  */
  assign n14394 = {n14393, cfg_cdiv};
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:191:58  */
  assign n14395 = {n14394, cfg_duty};
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:191:69  */
  assign n14396 = re_i ? n14395 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:200:16  */
  assign n14399 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:207:18  */
  assign n14401 = ~cfg_en;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:213:60  */
  assign n14406 = cnt_cdiv + 10'b0000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:210:9  */
  assign n14408 = cnt_tick ? 10'b0000000000 : n14406;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:209:7  */
  assign n14409 = n14449 ? n14408 : cnt_cdiv;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:207:7  */
  assign n14411 = n14401 ? 10'b0000000000 : n14409;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:218:18  */
  assign n14412 = ~cfg_en;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:221:58  */
  assign n14414 = cnt_duty + 8'b00000001;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:220:7  */
  assign n14415 = cnt_tick ? n14414 : cnt_duty;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:218:7  */
  assign n14417 = n14412 ? 8'b00000000 : n14415;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:225:18  */
  assign n14418 = ~cfg_en;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:225:48  */
  assign n14419 = $unsigned(cnt_duty) >= $unsigned(cfg_duty);
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:225:25  */
  assign n14420 = n14418 | n14419;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:225:7  */
  assign n14423 = n14420 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:235:34  */
  assign n14435 = cnt_cdiv == cfg_cdiv;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:235:19  */
  assign n14436 = n14435 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:180:5  */
  assign n14438 = we_i ? n14370 : cfg_en;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:180:5  */
  always @(posedge clk_i or posedge n14368)
    if (n14368)
      n14439 <= 1'b0;
    else
      n14439 <= n14438;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:180:5  */
  assign n14440 = we_i ? n14371 : cfg_prsc;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:180:5  */
  always @(posedge clk_i or posedge n14368)
    if (n14368)
      n14441 <= 3'b000;
    else
      n14441 <= n14440;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:180:5  */
  assign n14442 = we_i ? n14372 : cfg_cdiv;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:180:5  */
  always @(posedge clk_i or posedge n14368)
    if (n14368)
      n14443 <= 10'b0000000000;
    else
      n14443 <= n14442;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:180:5  */
  assign n14444 = we_i ? n14373 : cfg_duty;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:180:5  */
  always @(posedge clk_i or posedge n14368)
    if (n14368)
      n14445 <= 8'b00000000;
    else
      n14445 <= n14444;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:204:5  */
  always @(posedge clk_i or posedge n14399)
    if (n14399)
      n14446 <= 10'b0000000000;
    else
      n14446 <= n14411;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:204:5  */
  always @(posedge clk_i or posedge n14399)
    if (n14399)
      n14447 <= 8'b00000000;
    else
      n14447 <= n14417;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:204:5  */
  always @(posedge clk_i or posedge n14399)
    if (n14399)
      n14448 <= 1'b0;
    else
      n14448 <= n14423;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:209:23  */
  assign n14449 = clkgen_i[cfg_prsc * 1 +: 1]; //(Bmux)
endmodule

module neorv32_fifo_1_11_47ec8d98366433dc002e7721c9e37d5067547937
  (input  clk_i,
   input  rstn_i,
   input  clear_i,
   input  [10:0] wdata_i,
   input  we_i,
   input  re_i,
   output half_o,
   output free_o,
   output [10:0] rdata_o,
   output avail_o);
  wire [10:0] fifo_reg;
  wire we;
  wire re;
  wire match;
  wire empty;
  wire full;
  wire half;
  wire free;
  wire avail;
  wire w_pnt;
  wire w_nxt;
  wire r_pnt;
  wire r_nxt;
  wire n14304;
  wire n14305;
  wire n14307;
  wire n14308;
  wire n14310;
  wire n14320;
  wire n14322;
  wire n14323;
  wire n14325;
  wire n14327;
  wire n14328;
  wire n14330;
  wire n14331;
  wire n14333;
  wire n14334;
  wire n14335;
  wire n14342;
  wire [10:0] n14355;
  reg [10:0] n14356;
  reg n14357;
  reg n14358;
  reg n14361;
  reg n14362;
  reg n14363;
  assign half_o = n14361; //(module output)
  assign free_o = n14362; //(module output)
  assign rdata_o = fifo_reg; //(module output)
  assign avail_o = n14363; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:51:10  */
  assign fifo_reg = n14356; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:10  */
  assign we = n14307; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:14  */
  assign re = n14304; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:18  */
  assign match = n14331; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:25  */
  assign empty = match; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:32  */
  assign full = n14333; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:38  */
  assign half = full; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:44  */
  assign free = n14334; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:50  */
  assign avail = n14335; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:10  */
  assign w_pnt = n14357; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:17  */
  assign w_nxt = n14320; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:24  */
  assign r_pnt = n14358; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:31  */
  assign r_nxt = n14325; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:66:14  */
  assign n14304 = 1'b0 ? re_i : n14305;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:66:50  */
  assign n14305 = re_i & avail;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:67:14  */
  assign n14307 = 1'b0 ? we_i : n14308;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:67:50  */
  assign n14308 = we_i & free;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:74:16  */
  assign n14310 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:28  */
  assign n14320 = clear_i ? 1'b0 : n14323;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:88  */
  assign n14322 = w_pnt + 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:49  */
  assign n14323 = we ? n14322 : w_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:28  */
  assign n14325 = clear_i ? 1'b0 : n14328;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:88  */
  assign n14327 = r_pnt + 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:49  */
  assign n14328 = re ? n14327 : r_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:104:33  */
  assign n14330 = r_pnt == w_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:104:18  */
  assign n14331 = n14330 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:105:14  */
  assign n14333 = ~match;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:110:12  */
  assign n14334 = ~full;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:111:12  */
  assign n14335 = ~empty;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:242:18  */
  assign n14342 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:162:9  */
  assign n14355 = we ? wdata_i : fifo_reg;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:162:9  */
  always @(posedge clk_i)
    n14356 <= n14355;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:77:5  */
  always @(posedge clk_i or posedge n14310)
    if (n14310)
      n14357 <= 1'b0;
    else
      n14357 <= w_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:77:5  */
  always @(posedge clk_i or posedge n14310)
    if (n14310)
      n14358 <= 1'b0;
    else
      n14358 <= r_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14342)
    if (n14342)
      n14361 <= 1'b0;
    else
      n14361 <= half;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14342)
    if (n14342)
      n14362 <= 1'b0;
    else
      n14362 <= free;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14342)
    if (n14342)
      n14363 <= 1'b0;
    else
      n14363 <= avail;
endmodule

module neorv32_fifo_1_9_47ec8d98366433dc002e7721c9e37d5067547937
  (input  clk_i,
   input  rstn_i,
   input  clear_i,
   input  [8:0] wdata_i,
   input  we_i,
   input  re_i,
   output half_o,
   output free_o,
   output [8:0] rdata_o,
   output avail_o);
  wire [8:0] fifo_reg;
  wire we;
  wire re;
  wire match;
  wire empty;
  wire full;
  wire half;
  wire free;
  wire avail;
  wire w_pnt;
  wire w_nxt;
  wire r_pnt;
  wire r_nxt;
  wire n14239;
  wire n14240;
  wire n14242;
  wire n14243;
  wire n14245;
  wire n14255;
  wire n14257;
  wire n14258;
  wire n14260;
  wire n14262;
  wire n14263;
  wire n14265;
  wire n14266;
  wire n14268;
  wire n14269;
  wire n14270;
  wire n14277;
  wire [8:0] n14290;
  reg [8:0] n14291;
  reg n14292;
  reg n14293;
  reg n14296;
  reg n14297;
  reg n14298;
  assign half_o = n14296; //(module output)
  assign free_o = n14297; //(module output)
  assign rdata_o = fifo_reg; //(module output)
  assign avail_o = n14298; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:51:10  */
  assign fifo_reg = n14291; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:10  */
  assign we = n14242; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:14  */
  assign re = n14239; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:18  */
  assign match = n14266; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:25  */
  assign empty = match; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:32  */
  assign full = n14268; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:38  */
  assign half = full; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:44  */
  assign free = n14269; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:50  */
  assign avail = n14270; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:10  */
  assign w_pnt = n14292; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:17  */
  assign w_nxt = n14255; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:24  */
  assign r_pnt = n14293; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:31  */
  assign r_nxt = n14260; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:66:14  */
  assign n14239 = 1'b0 ? re_i : n14240;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:66:50  */
  assign n14240 = re_i & avail;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:67:14  */
  assign n14242 = 1'b0 ? we_i : n14243;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:67:50  */
  assign n14243 = we_i & free;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:74:16  */
  assign n14245 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:28  */
  assign n14255 = clear_i ? 1'b0 : n14258;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:88  */
  assign n14257 = w_pnt + 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:49  */
  assign n14258 = we ? n14257 : w_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:28  */
  assign n14260 = clear_i ? 1'b0 : n14263;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:88  */
  assign n14262 = r_pnt + 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:49  */
  assign n14263 = re ? n14262 : r_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:104:33  */
  assign n14265 = r_pnt == w_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:104:18  */
  assign n14266 = n14265 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:105:14  */
  assign n14268 = ~match;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:110:12  */
  assign n14269 = ~full;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:111:12  */
  assign n14270 = ~empty;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:242:18  */
  assign n14277 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:162:9  */
  assign n14290 = we ? wdata_i : fifo_reg;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:162:9  */
  always @(posedge clk_i)
    n14291 <= n14290;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:77:5  */
  always @(posedge clk_i or posedge n14245)
    if (n14245)
      n14292 <= 1'b0;
    else
      n14292 <= w_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:77:5  */
  always @(posedge clk_i or posedge n14245)
    if (n14245)
      n14293 <= 1'b0;
    else
      n14293 <= r_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14277)
    if (n14277)
      n14296 <= 1'b0;
    else
      n14296 <= half;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14277)
    if (n14277)
      n14297 <= 1'b0;
    else
      n14297 <= free;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14277)
    if (n14277)
      n14298 <= 1'b0;
    else
      n14298 <= avail;
endmodule

module neorv32_fifo_1_8_47ec8d98366433dc002e7721c9e37d5067547937
  (input  clk_i,
   input  rstn_i,
   input  clear_i,
   input  [7:0] wdata_i,
   input  we_i,
   input  re_i,
   output half_o,
   output free_o,
   output [7:0] rdata_o,
   output avail_o);
  wire [7:0] fifo_reg;
  wire we;
  wire re;
  wire match;
  wire empty;
  wire full;
  wire half;
  wire free;
  wire avail;
  wire w_pnt;
  wire w_nxt;
  wire r_pnt;
  wire r_nxt;
  wire n14174;
  wire n14175;
  wire n14177;
  wire n14178;
  wire n14180;
  wire n14190;
  wire n14192;
  wire n14193;
  wire n14195;
  wire n14197;
  wire n14198;
  wire n14200;
  wire n14201;
  wire n14203;
  wire n14204;
  wire n14205;
  wire n14212;
  wire [7:0] n14225;
  reg [7:0] n14226;
  reg n14227;
  reg n14228;
  reg n14231;
  reg n14232;
  reg n14233;
  assign half_o = n14231; //(module output)
  assign free_o = n14232; //(module output)
  assign rdata_o = fifo_reg; //(module output)
  assign avail_o = n14233; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:51:10  */
  assign fifo_reg = n14226; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:10  */
  assign we = n14177; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:14  */
  assign re = n14174; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:18  */
  assign match = n14201; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:25  */
  assign empty = match; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:32  */
  assign full = n14203; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:38  */
  assign half = full; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:44  */
  assign free = n14204; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:54:50  */
  assign avail = n14205; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:10  */
  assign w_pnt = n14227; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:17  */
  assign w_nxt = n14190; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:24  */
  assign r_pnt = n14228; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:57:31  */
  assign r_nxt = n14195; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:66:14  */
  assign n14174 = 1'b0 ? re_i : n14175;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:66:50  */
  assign n14175 = re_i & avail;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:67:14  */
  assign n14177 = 1'b0 ? we_i : n14178;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:67:50  */
  assign n14178 = we_i & free;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:74:16  */
  assign n14180 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:28  */
  assign n14190 = clear_i ? 1'b0 : n14193;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:88  */
  assign n14192 = w_pnt + 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:84:49  */
  assign n14193 = we ? n14192 : w_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:28  */
  assign n14195 = clear_i ? 1'b0 : n14198;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:88  */
  assign n14197 = r_pnt + 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:85:49  */
  assign n14198 = re ? n14197 : r_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:104:33  */
  assign n14200 = r_pnt == w_pnt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:104:18  */
  assign n14201 = n14200 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:105:14  */
  assign n14203 = ~match;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:110:12  */
  assign n14204 = ~full;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:111:12  */
  assign n14205 = ~empty;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:242:18  */
  assign n14212 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:162:9  */
  assign n14225 = we ? wdata_i : fifo_reg;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:162:9  */
  always @(posedge clk_i)
    n14226 <= n14225;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:77:5  */
  always @(posedge clk_i or posedge n14180)
    if (n14180)
      n14227 <= 1'b0;
    else
      n14227 <= w_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:77:5  */
  always @(posedge clk_i or posedge n14180)
    if (n14180)
      n14228 <= 1'b0;
    else
      n14228 <= r_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14212)
    if (n14212)
      n14231 <= 1'b0;
    else
      n14231 <= half;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14212)
    if (n14212)
      n14232 <= 1'b0;
    else
      n14232 <= free;
  /* ../../ext/neorv32/rtl/core/neorv32_fifo.vhd:246:7  */
  always @(posedge clk_i or posedge n14212)
    if (n14212)
      n14233 <= 1'b0;
    else
      n14233 <= avail;
endmodule

module neorv32_clint_swi
  (input  clk_i,
   input  rstn_i,
   input  en_i,
   input  rw_i,
   input  [31:0] wdata_i,
   output [31:0] rdata_o,
   output swi_o);
  wire rden_q;
  wire sip_q;
  wire n14150;
  wire n14152;
  wire n14153;
  wire n14163;
  reg n14165;
  wire n14166;
  reg n14167;
  wire [31:0] n14168;
  assign rdata_o = n14168; //(module output)
  assign swi_o = sip_q; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:427:10  */
  assign rden_q = n14165; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:427:18  */
  assign sip_q = n14167; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:435:16  */
  assign n14150 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:440:23  */
  assign n14152 = rw_i & en_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:441:25  */
  assign n14153 = wdata_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:448:23  */
  assign n14163 = rden_q ? sip_q : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:438:5  */
  always @(posedge clk_i or posedge n14150)
    if (n14150)
      n14165 <= 1'b0;
    else
      n14165 <= en_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:438:5  */
  assign n14166 = n14152 ? n14153 : sip_q;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:438:5  */
  always @(posedge clk_i or posedge n14150)
    if (n14150)
      n14167 <= 1'b0;
    else
      n14167 <= n14166;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:435:5  */
  assign n14168 = {31'b0000000000000000000000000000000, n14163};
endmodule

module neorv32_clint_mtimecmp
  (input  clk_i,
   input  rstn_i,
   input  en_i,
   input  rw_i,
   input  addr_i,
   input  [31:0] wdata_i,
   input  [63:0] mtime_i,
   output [31:0] rdata_o,
   output mti_o);
  wire [1:0] rden_q;
  wire [63:0] mtimecmp_q;
  wire cmp_lo_eq;
  wire cmp_lo_gt;
  wire cmp_lo_ge;
  wire cmp_hi_eq;
  wire cmp_hi_gt;
  wire n14077;
  wire n14079;
  wire n14080;
  wire n14081;
  wire n14082;
  wire n14083;
  wire [31:0] n14084;
  wire [31:0] n14085;
  wire [31:0] n14086;
  wire [31:0] n14087;
  wire [63:0] n14088;
  wire [1:0] n14090;
  wire [31:0] n14098;
  wire n14099;
  wire [31:0] n14100;
  wire [31:0] n14101;
  wire n14102;
  wire [31:0] n14103;
  wire n14106;
  wire n14108;
  wire n14109;
  wire n14110;
  wire [31:0] n14119;
  wire [31:0] n14120;
  wire n14121;
  wire n14122;
  wire [31:0] n14125;
  wire [31:0] n14126;
  wire n14127;
  wire n14128;
  wire [31:0] n14131;
  wire [31:0] n14132;
  wire n14133;
  wire n14134;
  wire [31:0] n14137;
  wire [31:0] n14138;
  wire n14139;
  wire n14140;
  reg [1:0] n14142;
  wire [63:0] n14143;
  reg [63:0] n14144;
  reg n14145;
  reg n14146;
  assign rdata_o = n14100; //(module output)
  assign mti_o = n14146; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:341:10  */
  assign rden_q = n14142; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:342:10  */
  assign mtimecmp_q = n14144; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:343:10  */
  assign cmp_lo_eq = n14122; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:343:21  */
  assign cmp_lo_gt = n14128; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:343:32  */
  assign cmp_lo_ge = n14145; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:343:43  */
  assign cmp_hi_eq = n14134; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:343:54  */
  assign cmp_hi_gt = n14140; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:351:16  */
  assign n14077 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:355:30  */
  assign n14079 = ~addr_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:355:25  */
  assign n14080 = en_i & n14079;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:356:25  */
  assign n14081 = en_i & addr_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:357:23  */
  assign n14082 = rw_i & en_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:358:20  */
  assign n14083 = ~addr_i;
  assign n14084 = mtimecmp_q[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:358:9  */
  assign n14085 = n14083 ? wdata_i : n14084;
  assign n14086 = mtimecmp_q[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:358:9  */
  assign n14087 = n14083 ? n14086 : wdata_i;
  assign n14088 = {n14087, n14085};
  assign n14090 = {n14081, n14080};
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:368:24  */
  assign n14098 = mtimecmp_q[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:368:51  */
  assign n14099 = rden_q[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:368:39  */
  assign n14100 = n14099 ? n14098 : n14103;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:369:24  */
  assign n14101 = mtimecmp_q[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:369:51  */
  assign n14102 = rden_q[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:368:62  */
  assign n14103 = n14102 ? n14101 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:377:16  */
  assign n14106 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:381:30  */
  assign n14108 = cmp_lo_gt | cmp_lo_eq;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:382:44  */
  assign n14109 = cmp_hi_eq & cmp_lo_ge;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:382:30  */
  assign n14110 = cmp_hi_gt | n14109;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:387:42  */
  assign n14119 = mtime_i[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:387:79  */
  assign n14120 = mtimecmp_q[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:387:58  */
  assign n14121 = n14119 == n14120;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:387:20  */
  assign n14122 = n14121 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:388:42  */
  assign n14125 = mtime_i[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:388:79  */
  assign n14126 = mtimecmp_q[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:388:58  */
  assign n14127 = $unsigned(n14125) > $unsigned(n14126);
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:388:20  */
  assign n14128 = n14127 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:389:42  */
  assign n14131 = mtime_i[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:389:79  */
  assign n14132 = mtimecmp_q[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:389:58  */
  assign n14133 = n14131 == n14132;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:389:20  */
  assign n14134 = n14133 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:390:42  */
  assign n14137 = mtime_i[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:390:79  */
  assign n14138 = mtimecmp_q[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:390:58  */
  assign n14139 = $unsigned(n14137) > $unsigned(n14138);
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:390:20  */
  assign n14140 = n14139 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:354:5  */
  always @(posedge clk_i or posedge n14077)
    if (n14077)
      n14142 <= 2'b00;
    else
      n14142 <= n14090;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:354:5  */
  assign n14143 = n14082 ? n14088 : mtimecmp_q;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:354:5  */
  always @(posedge clk_i or posedge n14077)
    if (n14077)
      n14144 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      n14144 <= n14143;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:380:5  */
  always @(posedge clk_i or posedge n14106)
    if (n14106)
      n14145 <= 1'b0;
    else
      n14145 <= n14108;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:380:5  */
  always @(posedge clk_i or posedge n14106)
    if (n14106)
      n14146 <= 1'b0;
    else
      n14146 <= n14110;
endmodule

module neorv32_clint_mtime
  (input  clk_i,
   input  rstn_i,
   input  en_i,
   input  rw_i,
   input  addr_i,
   input  [31:0] wdata_i,
   output [31:0] rdata_o,
   output [63:0] mtime_o);
  wire [1:0] re_q;
  wire [1:0] we_q;
  wire [31:0] mtime_lo_q;
  wire [31:0] mtime_hi_q;
  wire carry_q;
  wire [32:0] inc_lo;
  wire [32:0] inc_hi;
  wire n14020;
  wire n14022;
  wire n14023;
  wire n14024;
  wire n14025;
  wire n14026;
  wire n14027;
  wire n14028;
  wire n14029;
  wire n14030;
  wire [31:0] n14031;
  wire [31:0] n14032;
  wire n14033;
  wire n14034;
  wire [31:0] n14035;
  wire [31:0] n14036;
  wire [1:0] n14037;
  wire [1:0] n14039;
  wire [32:0] n14056;
  wire [32:0] n14058;
  wire [32:0] n14060;
  wire [32:0] n14061;
  wire [32:0] n14062;
  wire [63:0] n14063;
  wire n14064;
  wire [31:0] n14065;
  wire n14066;
  wire [31:0] n14067;
  reg [1:0] n14069;
  reg [1:0] n14070;
  reg [31:0] n14071;
  reg [31:0] n14072;
  reg n14073;
  assign rdata_o = n14065; //(module output)
  assign mtime_o = n14063; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:251:10  */
  assign re_q = n14069; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:252:10  */
  assign we_q = n14070; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:253:10  */
  assign mtime_lo_q = n14071; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:254:10  */
  assign mtime_hi_q = n14072; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:255:10  */
  assign carry_q = n14073; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:256:10  */
  assign inc_lo = n14058; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:257:10  */
  assign inc_hi = n14062; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:265:16  */
  assign n14020 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:272:23  */
  assign n14022 = en_i & rw_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:272:37  */
  assign n14023 = ~addr_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:272:32  */
  assign n14024 = n14022 & n14023;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:273:23  */
  assign n14025 = en_i & rw_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:273:32  */
  assign n14026 = n14025 & addr_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:274:28  */
  assign n14027 = ~addr_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:274:23  */
  assign n14028 = en_i & n14027;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:275:23  */
  assign n14029 = en_i & addr_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:277:15  */
  assign n14030 = we_q[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:280:29  */
  assign n14031 = inc_lo[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:277:7  */
  assign n14032 = n14030 ? wdata_i : n14031;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:282:27  */
  assign n14033 = inc_lo[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:284:15  */
  assign n14034 = we_q[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:287:29  */
  assign n14035 = inc_hi[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:284:7  */
  assign n14036 = n14034 ? wdata_i : n14035;
  assign n14037 = {n14029, n14028};
  assign n14039 = {n14026, n14024};
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:293:44  */
  assign n14056 = {1'b0, mtime_lo_q};
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:293:58  */
  assign n14058 = n14056 + 33'b000000000000000000000000000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:294:44  */
  assign n14060 = {1'b0, mtime_hi_q};
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:294:58  */
  assign n14061 = {32'b0, carry_q};  //  uext
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:294:58  */
  assign n14062 = n14060 + n14061;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:297:25  */
  assign n14063 = {mtime_hi_q, mtime_lo_q};
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:300:35  */
  assign n14064 = re_q[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:300:25  */
  assign n14065 = n14064 ? mtime_hi_q : n14067;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:301:35  */
  assign n14066 = re_q[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:300:46  */
  assign n14067 = n14066 ? mtime_lo_q : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:271:5  */
  always @(posedge clk_i or posedge n14020)
    if (n14020)
      n14069 <= 2'b00;
    else
      n14069 <= n14037;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:271:5  */
  always @(posedge clk_i or posedge n14020)
    if (n14020)
      n14070 <= 2'b00;
    else
      n14070 <= n14039;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:271:5  */
  always @(posedge clk_i or posedge n14020)
    if (n14020)
      n14071 <= 32'b00000000000000000000000000000000;
    else
      n14071 <= n14032;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:271:5  */
  always @(posedge clk_i or posedge n14020)
    if (n14020)
      n14072 <= 32'b00000000000000000000000000000000;
    else
      n14072 <= n14036;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:271:5  */
  always @(posedge clk_i or posedge n14020)
    if (n14020)
      n14073 <= 1'b0;
    else
      n14073 <= n14033;
endmodule

module neorv32_bus_reg_9159cb8bcee7fcb95582f140960cdae72788d326
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \host_req_i_host_req_i[addr] ,
   input  [31:0] \host_req_i_host_req_i[data] ,
   input  [3:0] \host_req_i_host_req_i[ben] ,
   input  \host_req_i_host_req_i[stb] ,
   input  \host_req_i_host_req_i[rw] ,
   input  \host_req_i_host_req_i[src] ,
   input  \host_req_i_host_req_i[priv] ,
   input  \host_req_i_host_req_i[amo] ,
   input  [3:0] \host_req_i_host_req_i[amoop] ,
   input  \host_req_i_host_req_i[fence] ,
   input  \host_req_i_host_req_i[sleep] ,
   input  \host_req_i_host_req_i[debug] ,
   input  [31:0] \device_rsp_i_device_rsp_i[data] ,
   input  \device_rsp_i_device_rsp_i[ack] ,
   input  \device_rsp_i_device_rsp_i[err] ,
   output [31:0] \host_rsp_o_host_rsp_o[data] ,
   output \host_rsp_o_host_rsp_o[ack] ,
   output \host_rsp_o_host_rsp_o[err] ,
   output [31:0] \device_req_o_device_req_o[addr] ,
   output [31:0] \device_req_o_device_req_o[data] ,
   output [3:0] \device_req_o_device_req_o[ben] ,
   output \device_req_o_device_req_o[stb] ,
   output \device_req_o_device_req_o[rw] ,
   output \device_req_o_device_req_o[src] ,
   output \device_req_o_device_req_o[priv] ,
   output \device_req_o_device_req_o[amo] ,
   output [3:0] \device_req_o_device_req_o[amoop] ,
   output \device_req_o_device_req_o[fence] ,
   output \device_req_o_device_req_o[sleep] ,
   output \device_req_o_device_req_o[debug] );
  wire [79:0] n13976;
  wire [31:0] n13978;
  wire n13979;
  wire n13980;
  wire [31:0] n13982;
  wire [31:0] n13983;
  wire [3:0] n13984;
  wire n13985;
  wire n13986;
  wire n13987;
  wire n13988;
  wire n13989;
  wire [3:0] n13990;
  wire n13991;
  wire n13992;
  wire n13993;
  wire [33:0] n13994;
  wire n13996;
  wire n13998;
  wire [79:0] n13999;
  wire n14000;
  wire [10:0] n14001;
  wire [67:0] n14002;
  wire [79:0] n14003;
  wire n14009;
  reg [33:0] n14015;
  reg [79:0] n14016;
  assign \host_rsp_o_host_rsp_o[data]  = n13978; //(module output)
  assign \host_rsp_o_host_rsp_o[ack]  = n13979; //(module output)
  assign \host_rsp_o_host_rsp_o[err]  = n13980; //(module output)
  assign \device_req_o_device_req_o[addr]  = n13982; //(module output)
  assign \device_req_o_device_req_o[data]  = n13983; //(module output)
  assign \device_req_o_device_req_o[ben]  = n13984; //(module output)
  assign \device_req_o_device_req_o[stb]  = n13985; //(module output)
  assign \device_req_o_device_req_o[rw]  = n13986; //(module output)
  assign \device_req_o_device_req_o[src]  = n13987; //(module output)
  assign \device_req_o_device_req_o[priv]  = n13988; //(module output)
  assign \device_req_o_device_req_o[amo]  = n13989; //(module output)
  assign \device_req_o_device_req_o[amoop]  = n13990; //(module output)
  assign \device_req_o_device_req_o[fence]  = n13991; //(module output)
  assign \device_req_o_device_req_o[sleep]  = n13992; //(module output)
  assign \device_req_o_device_req_o[debug]  = n13993; //(module output)
  assign n13976 = {\host_req_i_host_req_i[debug] , \host_req_i_host_req_i[sleep] , \host_req_i_host_req_i[fence] , \host_req_i_host_req_i[amoop] , \host_req_i_host_req_i[amo] , \host_req_i_host_req_i[priv] , \host_req_i_host_req_i[src] , \host_req_i_host_req_i[rw] , \host_req_i_host_req_i[stb] , \host_req_i_host_req_i[ben] , \host_req_i_host_req_i[data] , \host_req_i_host_req_i[addr] };
  assign n13978 = n14015[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1038:14  */
  assign n13979 = n14015[32]; // extract
  assign n13980 = n14015[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n13982 = n14016[31:0]; // extract
  assign n13983 = n14016[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n13984 = n14016[67:64]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:984:33  */
  assign n13985 = n14016[68]; // extract
  assign n13986 = n14016[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1038:14  */
  assign n13987 = n14016[70]; // extract
  assign n13988 = n14016[71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n13989 = n14016[72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n13990 = n14016[76:73]; // extract
  assign n13991 = n14016[77]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n13992 = n14016[78]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:920:33  */
  assign n13993 = n14016[79]; // extract
  assign n13994 = {\device_rsp_i_device_rsp_i[err] , \device_rsp_i_device_rsp_i[ack] , \device_rsp_i_device_rsp_i[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:252:18  */
  assign n13996 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:255:24  */
  assign n13998 = n13976[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:255:9  */
  assign n13999 = n13998 ? n13976 : n14016;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:258:40  */
  assign n14000 = n13976[68]; // extract
  assign n14001 = n13999[79:69]; // extract
  assign n14002 = n13999[67:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:847:3  */
  assign n14003 = {n14001, n14000, n14002};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:275:18  */
  assign n14009 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:277:7  */
  always @(posedge clk_i or posedge n14009)
    if (n14009)
      n14015 <= 34'b0000000000000000000000000000000000;
    else
      n14015 <= n13994;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:254:7  */
  always @(posedge clk_i or posedge n13996)
    if (n13996)
      n14016 <= 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      n14016 <= n14003;
endmodule

module neorv32_bus_reg_1489f923c4dca729178b3e3233458550d8dddf29
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \host_req_i_host_req_i[addr] ,
   input  [31:0] \host_req_i_host_req_i[data] ,
   input  [3:0] \host_req_i_host_req_i[ben] ,
   input  \host_req_i_host_req_i[stb] ,
   input  \host_req_i_host_req_i[rw] ,
   input  \host_req_i_host_req_i[src] ,
   input  \host_req_i_host_req_i[priv] ,
   input  \host_req_i_host_req_i[amo] ,
   input  [3:0] \host_req_i_host_req_i[amoop] ,
   input  \host_req_i_host_req_i[fence] ,
   input  \host_req_i_host_req_i[sleep] ,
   input  \host_req_i_host_req_i[debug] ,
   input  [31:0] \device_rsp_i_device_rsp_i[data] ,
   input  \device_rsp_i_device_rsp_i[ack] ,
   input  \device_rsp_i_device_rsp_i[err] ,
   output [31:0] \host_rsp_o_host_rsp_o[data] ,
   output \host_rsp_o_host_rsp_o[ack] ,
   output \host_rsp_o_host_rsp_o[err] ,
   output [31:0] \device_req_o_device_req_o[addr] ,
   output [31:0] \device_req_o_device_req_o[data] ,
   output [3:0] \device_req_o_device_req_o[ben] ,
   output \device_req_o_device_req_o[stb] ,
   output \device_req_o_device_req_o[rw] ,
   output \device_req_o_device_req_o[src] ,
   output \device_req_o_device_req_o[priv] ,
   output \device_req_o_device_req_o[amo] ,
   output [3:0] \device_req_o_device_req_o[amoop] ,
   output \device_req_o_device_req_o[fence] ,
   output \device_req_o_device_req_o[sleep] ,
   output \device_req_o_device_req_o[debug] );
  wire [79:0] n13957;
  wire [31:0] n13959;
  wire n13960;
  wire n13961;
  wire [31:0] n13963;
  wire [31:0] n13964;
  wire [3:0] n13965;
  wire n13966;
  wire n13967;
  wire n13968;
  wire n13969;
  wire n13970;
  wire [3:0] n13971;
  wire n13972;
  wire n13973;
  wire n13974;
  wire [33:0] n13975;
  assign \host_rsp_o_host_rsp_o[data]  = n13959; //(module output)
  assign \host_rsp_o_host_rsp_o[ack]  = n13960; //(module output)
  assign \host_rsp_o_host_rsp_o[err]  = n13961; //(module output)
  assign \device_req_o_device_req_o[addr]  = n13963; //(module output)
  assign \device_req_o_device_req_o[data]  = n13964; //(module output)
  assign \device_req_o_device_req_o[ben]  = n13965; //(module output)
  assign \device_req_o_device_req_o[stb]  = n13966; //(module output)
  assign \device_req_o_device_req_o[rw]  = n13967; //(module output)
  assign \device_req_o_device_req_o[src]  = n13968; //(module output)
  assign \device_req_o_device_req_o[priv]  = n13969; //(module output)
  assign \device_req_o_device_req_o[amo]  = n13970; //(module output)
  assign \device_req_o_device_req_o[amoop]  = n13971; //(module output)
  assign \device_req_o_device_req_o[fence]  = n13972; //(module output)
  assign \device_req_o_device_req_o[sleep]  = n13973; //(module output)
  assign \device_req_o_device_req_o[debug]  = n13974; //(module output)
  assign n13957 = {\host_req_i_host_req_i[debug] , \host_req_i_host_req_i[sleep] , \host_req_i_host_req_i[fence] , \host_req_i_host_req_i[amoop] , \host_req_i_host_req_i[amo] , \host_req_i_host_req_i[priv] , \host_req_i_host_req_i[src] , \host_req_i_host_req_i[rw] , \host_req_i_host_req_i[stb] , \host_req_i_host_req_i[ben] , \host_req_i_host_req_i[data] , \host_req_i_host_req_i[addr] };
  assign n13959 = n13975[31:0]; // extract
  assign n13960 = n13975[32]; // extract
  assign n13961 = n13975[33]; // extract
  assign n13963 = n13957[31:0]; // extract
  assign n13964 = n13957[63:32]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:837:5  */
  assign n13965 = n13957[67:64]; // extract
  assign n13966 = n13957[68]; // extract
  assign n13967 = n13957[69]; // extract
  assign n13968 = n13957[70]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  assign n13969 = n13957[71]; // extract
  assign n13970 = n13957[72]; // extract
  assign n13971 = n13957[76:73]; // extract
  assign n13972 = n13957[77]; // extract
  assign n13973 = n13957[78]; // extract
  assign n13974 = n13957[79]; // extract
  assign n13975 = {\device_rsp_i_device_rsp_i[err] , \device_rsp_i_device_rsp_i[ack] , \device_rsp_i_device_rsp_i[data] };
endmodule

module neorv32_cache_bus_16_64_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  rstn_i,
   input  clk_i,
   input  [31:0] \host_req_i_host_req_i[addr] ,
   input  [31:0] \host_req_i_host_req_i[data] ,
   input  [3:0] \host_req_i_host_req_i[ben] ,
   input  \host_req_i_host_req_i[stb] ,
   input  \host_req_i_host_req_i[rw] ,
   input  \host_req_i_host_req_i[src] ,
   input  \host_req_i_host_req_i[priv] ,
   input  \host_req_i_host_req_i[amo] ,
   input  [3:0] \host_req_i_host_req_i[amoop] ,
   input  \host_req_i_host_req_i[fence] ,
   input  \host_req_i_host_req_i[sleep] ,
   input  \host_req_i_host_req_i[debug] ,
   input  [31:0] \bus_rsp_i_bus_rsp_i[data] ,
   input  \bus_rsp_i_bus_rsp_i[ack] ,
   input  \bus_rsp_i_bus_rsp_i[err] ,
   input  cmd_sync_i,
   input  cmd_miss_i,
   input  dirty_i,
   input  [31:0] base_i,
   input  [31:0] rdata_i,
   output [31:0] \bus_req_o_bus_req_o[addr] ,
   output [31:0] \bus_req_o_bus_req_o[data] ,
   output [3:0] \bus_req_o_bus_req_o[ben] ,
   output \bus_req_o_bus_req_o[stb] ,
   output \bus_req_o_bus_req_o[rw] ,
   output \bus_req_o_bus_req_o[src] ,
   output \bus_req_o_bus_req_o[priv] ,
   output \bus_req_o_bus_req_o[amo] ,
   output [3:0] \bus_req_o_bus_req_o[amoop] ,
   output \bus_req_o_bus_req_o[fence] ,
   output \bus_req_o_bus_req_o[sleep] ,
   output \bus_req_o_bus_req_o[debug] ,
   output cmd_busy_o,
   output inval_o,
   output new_o,
   output [31:0] addr_o,
   output [3:0] we_o,
   output swe_o,
   output [31:0] wdata_o,
   output wstat_o);
  wire [79:0] n13728;
  wire [31:0] n13730;
  wire [31:0] n13731;
  wire [3:0] n13732;
  wire n13733;
  wire n13734;
  wire n13735;
  wire n13736;
  wire n13737;
  wire [3:0] n13738;
  wire n13739;
  wire n13740;
  wire n13741;
  wire [33:0] n13742;
  wire [3:0] state;
  wire [3:0] state_nxt;
  wire [29:0] haddr;
  wire [29:0] baddr;
  wire [29:0] addr;
  wire [29:0] addr_nxt;
  wire [21:0] n13751;
  wire [21:0] n13754;
  wire [3:0] n13755;
  wire n13758;
  wire [29:0] n13770;
  wire [21:0] n13774;
  wire [3:0] n13775;
  wire [25:0] n13776;
  wire [3:0] n13777;
  wire [29:0] n13778;
  wire [31:0] n13780;
  wire [31:0] n13781;
  wire n13782;
  wire [21:0] n13783;
  wire [3:0] n13784;
  wire [25:0] n13785;
  wire [3:0] n13786;
  wire [29:0] n13787;
  wire [31:0] n13789;
  localparam [79:0] n13790 = 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire n13804;
  wire n13807;
  wire n13808;
  wire n13810;
  wire n13811;
  wire [3:0] n13814;
  wire [3:0] n13816;
  wire n13818;
  wire [3:0] n13819;
  wire [21:0] n13820;
  wire n13822;
  wire n13826;
  wire n13828;
  wire n13829;
  wire n13830;
  wire [3:0] n13831;
  wire [3:0] n13833;
  wire n13841;
  wire n13843;
  wire n13845;
  wire n13846;
  wire n13847;
  wire n13848;
  wire n13849;
  wire n13850;
  wire [3:0] n13853;
  wire [3:0] n13854;
  wire [3:0] n13855;
  wire [3:0] n13856;
  wire n13858;
  wire n13860;
  wire n13862;
  wire n13864;
  wire n13869;
  wire n13871;
  wire [21:0] n13872;
  wire [3:0] n13873;
  wire [3:0] n13875;
  wire n13883;
  wire n13885;
  wire n13887;
  wire n13888;
  wire n13889;
  wire n13890;
  wire n13891;
  wire n13892;
  wire n13895;
  wire [3:0] n13898;
  wire n13900;
  wire [9:0] n13901;
  wire n13902;
  reg n13903;
  wire n13904;
  reg n13905;
  reg n13906;
  reg n13910;
  reg n13914;
  reg [3:0] n13918;
  reg n13922;
  reg [3:0] n13932;
  wire [21:0] n13936;
  reg [21:0] n13937;
  wire [3:0] n13938;
  reg [3:0] n13939;
  wire [3:0] n13940;
  reg [3:0] n13941;
  wire n13947;
  wire n13948;
  reg [3:0] n13950;
  wire [29:0] n13952;
  wire [29:0] n13953;
  reg [29:0] n13954;
  wire [29:0] n13955;
  wire [79:0] n13956;
  assign \bus_req_o_bus_req_o[addr]  = n13730; //(module output)
  assign \bus_req_o_bus_req_o[data]  = n13731; //(module output)
  assign \bus_req_o_bus_req_o[ben]  = n13732; //(module output)
  assign \bus_req_o_bus_req_o[stb]  = n13733; //(module output)
  assign \bus_req_o_bus_req_o[rw]  = n13734; //(module output)
  assign \bus_req_o_bus_req_o[src]  = n13735; //(module output)
  assign \bus_req_o_bus_req_o[priv]  = n13736; //(module output)
  assign \bus_req_o_bus_req_o[amo]  = n13737; //(module output)
  assign \bus_req_o_bus_req_o[amoop]  = n13738; //(module output)
  assign \bus_req_o_bus_req_o[fence]  = n13739; //(module output)
  assign \bus_req_o_bus_req_o[sleep]  = n13740; //(module output)
  assign \bus_req_o_bus_req_o[debug]  = n13741; //(module output)
  assign cmd_busy_o = n13948; //(module output)
  assign inval_o = n13910; //(module output)
  assign new_o = n13914; //(module output)
  assign addr_o = n13780; //(module output)
  assign we_o = n13918; //(module output)
  assign swe_o = n13922; //(module output)
  assign wdata_o = n13781; //(module output)
  assign wstat_o = n13782; //(module output)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:670:33  */
  assign n13728 = {\host_req_i_host_req_i[debug] , \host_req_i_host_req_i[sleep] , \host_req_i_host_req_i[fence] , \host_req_i_host_req_i[amoop] , \host_req_i_host_req_i[amo] , \host_req_i_host_req_i[priv] , \host_req_i_host_req_i[src] , \host_req_i_host_req_i[rw] , \host_req_i_host_req_i[stb] , \host_req_i_host_req_i[ben] , \host_req_i_host_req_i[data] , \host_req_i_host_req_i[addr] };
  assign n13730 = n13956[31:0]; // extract
  assign n13731 = n13956[63:32]; // extract
  assign n13732 = n13956[67:64]; // extract
  assign n13733 = n13956[68]; // extract
  assign n13734 = n13956[69]; // extract
  assign n13735 = n13956[70]; // extract
  assign n13736 = n13956[71]; // extract
  assign n13737 = n13956[72]; // extract
  assign n13738 = n13956[76:73]; // extract
  assign n13739 = n13956[77]; // extract
  assign n13740 = n13956[78]; // extract
  assign n13741 = n13956[79]; // extract
  assign n13742 = {\bus_rsp_i_bus_rsp_i[err] , \bus_rsp_i_bus_rsp_i[ack] , \bus_rsp_i_bus_rsp_i[data] };
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:802:10  */
  assign state = n13950; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:802:24  */
  assign state_nxt = n13932; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:810:10  */
  assign haddr = n13952; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:810:17  */
  assign baddr = n13953; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:810:24  */
  assign addr = n13954; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:810:30  */
  assign addr_nxt = n13955; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:817:31  */
  assign n13751 = n13728[31:10]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:822:22  */
  assign n13754 = base_i[31:10]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:823:22  */
  assign n13755 = base_i[9:6]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:831:16  */
  assign n13758 = ~rstn_i;
  assign n13770 = {4'b0000, 4'b0000, 22'b0000000000000000000000};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:855:21  */
  assign n13774 = addr[21:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:855:32  */
  assign n13775 = addr[25:22]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:855:25  */
  assign n13776 = {n13774, n13775};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:855:43  */
  assign n13777 = addr[29:26]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:855:36  */
  assign n13778 = {n13776, n13777};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:855:47  */
  assign n13780 = {n13778, 2'b00};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:858:26  */
  assign n13781 = n13742[31:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:859:26  */
  assign n13782 = n13742[33]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:867:29  */
  assign n13783 = addr[21:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:867:40  */
  assign n13784 = addr[25:22]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:867:33  */
  assign n13785 = {n13783, n13784};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:867:51  */
  assign n13786 = addr[29:26]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:867:44  */
  assign n13787 = {n13785, n13786};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:867:55  */
  assign n13789 = {n13787, 2'b00};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:874:35  */
  assign n13804 = n13728[79]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:875:15  */
  assign n13807 = state == 4'b0000;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:876:37  */
  assign n13808 = n13728[78]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:875:5  */
  assign n13810 = n13807 ? n13808 : 1'b0;
  assign n13811 = n13790[77]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:889:9  */
  assign n13814 = cmd_miss_i ? 4'b0001 : state;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:887:9  */
  assign n13816 = cmd_sync_i ? 4'b0111 : n13814;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:884:7  */
  assign n13818 = state == 4'b0000;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:896:31  */
  assign n13819 = baddr[25:22]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:901:33  */
  assign n13820 = haddr[21:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:893:7  */
  assign n13822 = state == 4'b0001;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:906:7  */
  assign n13826 = state == 4'b0010;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:918:23  */
  assign n13828 = n13742[32]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:918:48  */
  assign n13829 = n13742[33]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:918:34  */
  assign n13830 = n13828 | n13829;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:919:59  */
  assign n13831 = addr[29:26]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:919:64  */
  assign n13833 = n13831 + 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n13841 = addr[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n13843 = 1'b1 & n13841;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n13845 = addr[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n13846 = n13843 & n13845;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n13847 = addr[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n13848 = n13846 & n13847;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n13849 = addr[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n13850 = n13848 & n13849;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:920:11  */
  assign n13853 = n13850 ? 4'b0000 : 4'b0010;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:918:9  */
  assign n13854 = n13830 ? n13853 : state;
  assign n13855 = addr[29:26]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:918:9  */
  assign n13856 = n13830 ? n13833 : n13855;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:912:7  */
  assign n13858 = state == 4'b0011;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:928:7  */
  assign n13860 = state == 4'b0100;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:937:7  */
  assign n13862 = state == 4'b0101;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:947:7  */
  assign n13864 = state == 4'b0110;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:965:7  */
  assign n13869 = state == 4'b0111;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:972:7  */
  assign n13871 = state == 4'b1000;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:978:31  */
  assign n13872 = baddr[21:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:983:59  */
  assign n13873 = addr[25:22]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:983:64  */
  assign n13875 = n13873 + 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n13883 = addr[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n13885 = 1'b1 & n13883;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n13887 = addr[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n13888 = n13885 & n13887;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n13889 = addr[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n13890 = n13888 & n13889;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n13891 = addr[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n13892 = n13890 & n13891;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:984:11  */
  assign n13895 = n13892 ? 1'b0 : n13811;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:984:11  */
  assign n13898 = n13892 ? 4'b0000 : 4'b1000;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:976:7  */
  assign n13900 = state == 4'b1001;
  assign n13901 = {n13900, n13871, n13869, n13864, n13862, n13860, n13858, n13826, n13822, n13818};
  assign n13902 = n13790[68]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13903 = n13902;
      10'b0100000000: n13903 = n13902;
      10'b0010000000: n13903 = n13902;
      10'b0001000000: n13903 = n13902;
      10'b0000100000: n13903 = n13902;
      10'b0000010000: n13903 = n13902;
      10'b0000001000: n13903 = n13902;
      10'b0000000100: n13903 = 1'b1;
      10'b0000000010: n13903 = n13902;
      10'b0000000001: n13903 = n13902;
      default: n13903 = n13902;
    endcase
  assign n13904 = n13790[69]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13905 = n13904;
      10'b0100000000: n13905 = n13904;
      10'b0010000000: n13905 = n13904;
      10'b0001000000: n13905 = n13904;
      10'b0000100000: n13905 = n13904;
      10'b0000010000: n13905 = n13904;
      10'b0000001000: n13905 = 1'b0;
      10'b0000000100: n13905 = 1'b0;
      10'b0000000010: n13905 = n13904;
      10'b0000000001: n13905 = n13904;
      default: n13905 = n13904;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13906 = n13895;
      10'b0100000000: n13906 = n13811;
      10'b0010000000: n13906 = 1'b1;
      10'b0001000000: n13906 = n13811;
      10'b0000100000: n13906 = n13811;
      10'b0000010000: n13906 = n13811;
      10'b0000001000: n13906 = n13811;
      10'b0000000100: n13906 = n13811;
      10'b0000000010: n13906 = n13811;
      10'b0000000001: n13906 = n13811;
      default: n13906 = n13811;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13910 = 1'b1;
      10'b0100000000: n13910 = 1'b0;
      10'b0010000000: n13910 = 1'b0;
      10'b0001000000: n13910 = 1'b0;
      10'b0000100000: n13910 = 1'b0;
      10'b0000010000: n13910 = 1'b0;
      10'b0000001000: n13910 = 1'b0;
      10'b0000000100: n13910 = 1'b0;
      10'b0000000010: n13910 = 1'b0;
      10'b0000000001: n13910 = 1'b0;
      default: n13910 = 1'b0;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13914 = 1'b0;
      10'b0100000000: n13914 = 1'b0;
      10'b0010000000: n13914 = 1'b0;
      10'b0001000000: n13914 = 1'b0;
      10'b0000100000: n13914 = 1'b0;
      10'b0000010000: n13914 = 1'b0;
      10'b0000001000: n13914 = 1'b1;
      10'b0000000100: n13914 = 1'b0;
      10'b0000000010: n13914 = 1'b0;
      10'b0000000001: n13914 = 1'b0;
      default: n13914 = 1'b0;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13918 = 4'b0000;
      10'b0100000000: n13918 = 4'b0000;
      10'b0010000000: n13918 = 4'b0000;
      10'b0001000000: n13918 = 4'b0000;
      10'b0000100000: n13918 = 4'b0000;
      10'b0000010000: n13918 = 4'b0000;
      10'b0000001000: n13918 = 4'b1111;
      10'b0000000100: n13918 = 4'b0000;
      10'b0000000010: n13918 = 4'b0000;
      10'b0000000001: n13918 = 4'b0000;
      default: n13918 = 4'b0000;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13922 = 1'b0;
      10'b0100000000: n13922 = 1'b0;
      10'b0010000000: n13922 = 1'b0;
      10'b0001000000: n13922 = 1'b0;
      10'b0000100000: n13922 = 1'b0;
      10'b0000010000: n13922 = 1'b0;
      10'b0000001000: n13922 = 1'b1;
      10'b0000000100: n13922 = 1'b0;
      10'b0000000010: n13922 = 1'b0;
      10'b0000000001: n13922 = 1'b0;
      default: n13922 = 1'b0;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13932 = n13898;
      10'b0100000000: n13932 = 4'b1001;
      10'b0010000000: n13932 = 4'b1000;
      10'b0001000000: n13932 = 4'b0000;
      10'b0000100000: n13932 = 4'b0000;
      10'b0000010000: n13932 = 4'b0000;
      10'b0000001000: n13932 = n13854;
      10'b0000000100: n13932 = 4'b0011;
      10'b0000000010: n13932 = 4'b0010;
      10'b0000000001: n13932 = n13816;
      default: n13932 = 4'b0000;
    endcase
  assign n13936 = addr[21:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13937 = n13872;
      10'b0100000000: n13937 = n13936;
      10'b0010000000: n13937 = n13936;
      10'b0001000000: n13937 = n13936;
      10'b0000100000: n13937 = n13936;
      10'b0000010000: n13937 = n13936;
      10'b0000001000: n13937 = n13936;
      10'b0000000100: n13937 = n13936;
      10'b0000000010: n13937 = n13820;
      10'b0000000001: n13937 = n13936;
      default: n13937 = n13936;
    endcase
  assign n13938 = addr[25:22]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13939 = n13875;
      10'b0100000000: n13939 = n13938;
      10'b0010000000: n13939 = 4'b0000;
      10'b0001000000: n13939 = n13938;
      10'b0000100000: n13939 = n13938;
      10'b0000010000: n13939 = n13938;
      10'b0000001000: n13939 = n13938;
      10'b0000000100: n13939 = n13938;
      10'b0000000010: n13939 = n13819;
      10'b0000000001: n13939 = n13938;
      default: n13939 = n13938;
    endcase
  assign n13940 = addr[29:26]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:882:5  */
  always @*
    case (n13901)
      10'b1000000000: n13941 = n13940;
      10'b0100000000: n13941 = n13940;
      10'b0010000000: n13941 = n13940;
      10'b0001000000: n13941 = n13940;
      10'b0000100000: n13941 = n13940;
      10'b0000010000: n13941 = n13940;
      10'b0000001000: n13941 = n13856;
      10'b0000000100: n13941 = n13940;
      10'b0000000010: n13941 = n13940;
      10'b0000000001: n13941 = 4'b0000;
      default: n13941 = n13940;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:1001:33  */
  assign n13947 = state == 4'b0000;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:1001:21  */
  assign n13948 = n13947 ? 1'b0 : 1'b1;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:837:5  */
  always @(posedge clk_i or posedge n13758)
    if (n13758)
      n13950 <= 4'b0000;
    else
      n13950 <= state_nxt;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:831:5  */
  assign n13952 = {4'b0000, 4'b0000, n13751};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:831:5  */
  assign n13953 = {4'b0000, n13755, n13754};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:837:5  */
  always @(posedge clk_i or posedge n13758)
    if (n13758)
      n13954 <= n13770;
    else
      n13954 <= addr_nxt;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:831:5  */
  assign n13955 = {n13941, n13939, n13937};
  assign n13956 = {n13804, n13810, n13906, 4'b0000, 1'b0, 1'b0, 1'b0, n13905, n13903, 4'b1111, rdata_i, n13789};
endmodule

module neorv32_cache_memory_16_64_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  rstn_i,
   input  clk_i,
   input  inval_i,
   input  new_i,
   input  dirty_i,
   input  [31:0] addr_i,
   input  [3:0] we_i,
   input  swe_i,
   input  [31:0] wdata_i,
   input  wstat_i,
   output hit_o,
   output dirty_o,
   output [31:0] base_o,
   output [31:0] rdata_o,
   output rstat_o);
  wire [15:0] valid_mem;
  wire valid_mem_rd;
  wire [21:0] tag_mem_rd;
  wire [31:0] data_mem_rd;
  wire stat_mem_rd;
  wire [21:0] acc_tag;
  wire [21:0] acc_tag_ff;
  wire [3:0] acc_idx;
  wire [3:0] acc_idx_ff;
  wire [3:0] acc_off;
  wire [7:0] acc_adr;
  wire mem_wen;
  wire [47:0] mem_bm;
  wire [47:0] mem_dout;
  wire [7:0] mem_addr;
  wire [21:0] n13445;
  wire [3:0] n13446;
  wire [3:0] n13447;
  wire [7:0] n13448;
  wire n13450;
  wire n13460;
  wire [15:0] n13474;
  wire [15:0] n13480;
  wire n13516;
  wire n13517;
  wire n13518;
  wire n13523;
  localparam n13526 = 1'b1;
  localparam n13527 = 1'b1;
  wire [15:0] n13529;
  wire [47:0] n13530;
  localparam n13531 = 1'b1;
  localparam n13533 = 1'b0;
  localparam n13534 = 1'b0;
  localparam n13535 = 1'b0;
  localparam n13536 = 1'b0;
  localparam n13537 = 1'b0;
  localparam [7:0] n13538 = 8'b00000000;
  localparam [47:0] n13539 = 48'b000000000000000000000000000000000000000000000000;
  localparam [47:0] n13540 = 48'b000000000000000000000000000000000000000000000000;
  wire n13544;
  wire n13545;
  wire n13548;
  wire n13549;
  wire [7:0] n13550;
  wire n13553;
  wire n13554;
  wire [7:0] n13555;
  wire n13558;
  wire n13559;
  wire [7:0] n13560;
  wire n13563;
  wire n13564;
  wire [7:0] n13565;
  wire [31:0] n13568;
  wire n13569;
  wire n13570;
  reg [15:0] n13571;
  wire n13573;
  wire n13574;
  reg n13575;
  reg [21:0] n13582;
  reg [3:0] n13583;
  wire [47:0] n13584;
  wire [31:0] n13585;
  reg [21:0] n13587; // mem_rd
  wire n13589;
  wire n13590;
  wire n13591;
  wire n13592;
  wire n13593;
  wire n13594;
  wire n13595;
  wire n13596;
  wire n13597;
  wire n13598;
  wire n13599;
  wire n13600;
  wire n13601;
  wire n13602;
  wire n13603;
  wire n13604;
  wire n13605;
  wire n13606;
  wire n13607;
  wire n13608;
  wire n13609;
  wire n13610;
  wire n13611;
  wire n13612;
  wire n13613;
  wire n13614;
  wire n13615;
  wire n13616;
  wire n13617;
  wire n13618;
  wire n13619;
  wire n13620;
  wire n13621;
  wire n13622;
  wire n13623;
  wire n13624;
  wire n13625;
  wire n13626;
  wire n13627;
  wire n13628;
  wire n13629;
  wire n13630;
  wire n13631;
  wire n13632;
  wire n13633;
  wire n13634;
  wire n13635;
  wire n13636;
  wire n13637;
  wire n13638;
  wire n13639;
  wire n13640;
  wire n13641;
  wire n13642;
  wire n13643;
  wire n13644;
  wire n13645;
  wire n13646;
  wire n13647;
  wire n13648;
  wire n13649;
  wire n13650;
  wire n13651;
  wire n13652;
  wire n13653;
  wire n13654;
  wire n13655;
  wire n13656;
  wire [15:0] n13657;
  wire n13658;
  wire n13659;
  wire n13660;
  wire n13661;
  wire n13662;
  wire n13663;
  wire n13664;
  wire n13665;
  wire n13666;
  wire n13667;
  wire n13668;
  wire n13669;
  wire n13670;
  wire n13671;
  wire n13672;
  wire n13673;
  wire n13674;
  wire n13675;
  wire n13676;
  wire n13677;
  wire n13678;
  wire n13679;
  wire n13680;
  wire n13681;
  wire n13682;
  wire n13683;
  wire n13684;
  wire n13685;
  wire n13686;
  wire n13687;
  wire n13688;
  wire n13689;
  wire n13690;
  wire n13691;
  wire n13692;
  wire n13693;
  wire n13694;
  wire n13695;
  wire n13696;
  wire n13697;
  wire n13698;
  wire n13699;
  wire n13700;
  wire n13701;
  wire n13702;
  wire n13703;
  wire n13704;
  wire n13705;
  wire n13706;
  wire n13707;
  wire n13708;
  wire n13709;
  wire n13710;
  wire n13711;
  wire n13712;
  wire n13713;
  wire n13714;
  wire n13715;
  wire n13716;
  wire n13717;
  wire n13718;
  wire n13719;
  wire n13720;
  wire n13721;
  wire n13722;
  wire n13723;
  wire n13724;
  wire n13725;
  wire [15:0] n13726;
  wire n13727;
  assign hit_o = n13518; //(module output)
  assign dirty_o = n13523; //(module output)
  assign base_o = n13585; //(module output)
  assign rdata_o = data_mem_rd; //(module output)
  assign rstat_o = n13570; //(module output)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:579:10  */
  assign valid_mem = n13571; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:580:10  */
  assign valid_mem_rd = n13575; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:585:10  */
  assign tag_mem_rd = n13587; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:588:10  */
  assign data_mem_rd = n13568; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:591:10  */
  assign stat_mem_rd = n13569; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:594:10  */
  assign acc_tag = n13445; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:594:19  */
  assign acc_tag_ff = n13582; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:595:10  */
  assign acc_idx = n13446; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:595:19  */
  assign acc_idx_ff = n13583; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:596:10  */
  assign acc_off = n13447; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:722:50  */
  assign acc_adr = n13448; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:621:10  */
  assign mem_wen = n13545; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:622:10  */
  assign mem_bm = n13584; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:624:10  */
  assign mem_addr = acc_adr; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:632:20  */
  assign n13445 = addr_i[31:10]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:633:20  */
  assign n13446 = addr_i[9:6]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:634:20  */
  assign n13447 = addr_i[5:2]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:635:22  */
  assign n13448 = {acc_idx, acc_off};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:640:16  */
  assign n13450 = ~rstn_i;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:654:16  */
  assign n13460 = ~rstn_i;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:662:9  */
  assign n13474 = inval_i ? n13726 : valid_mem;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:658:7  */
  assign n13480 = new_i ? n13657 : n13474;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:691:60  */
  assign n13516 = tag_mem_rd == acc_tag_ff;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:691:44  */
  assign n13517 = n13516 & valid_mem_rd;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:691:18  */
  assign n13518 = n13517 ? 1'b1 : 1'b0;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:692:18  */
  assign n13523 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:702:3  */
  RM_IHPSG13_1P_256x48_c2_bm_bist mem (
    .A_CLK(clk_i),
    .A_MEN(n13526),
    .A_WEN(mem_wen),
    .A_REN(n13527),
    .A_ADDR(mem_addr),
    .A_DIN(n13530),
    .A_DLY(n13531),
    .A_BM(mem_bm),
    .A_BIST_CLK(n13533),
    .A_BIST_EN(n13534),
    .A_BIST_MEN(n13535),
    .A_BIST_WEN(n13536),
    .A_BIST_REN(n13537),
    .A_BIST_ADDR(n13538),
    .A_BIST_DIN(n13539),
    .A_BIST_BM(n13540),
    .A_DOUT(mem_dout));
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:709:31  */
  assign n13529 = {15'b000000000000000, wstat_i};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:709:41  */
  assign n13530 = {n13529, wdata_i};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:723:28  */
  assign n13544 = we_i == 4'b0000;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:723:18  */
  assign n13545 = n13544 ? 1'b0 : 1'b1;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:724:40  */
  assign n13548 = we_i[0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:724:44  */
  assign n13549 = ~n13548;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:724:31  */
  assign n13550 = n13549 ? 8'b00000000 : 8'b11111111;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:725:41  */
  assign n13553 = we_i[1]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:725:45  */
  assign n13554 = ~n13553;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:725:32  */
  assign n13555 = n13554 ? 8'b00000000 : 8'b11111111;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:726:42  */
  assign n13558 = we_i[2]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:726:46  */
  assign n13559 = ~n13558;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:726:33  */
  assign n13560 = n13559 ? 8'b00000000 : 8'b11111111;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:727:42  */
  assign n13563 = we_i[3]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:727:46  */
  assign n13564 = ~n13563;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:727:33  */
  assign n13565 = n13564 ? 8'b00000000 : 8'b11111111;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:730:26  */
  assign n13568 = mem_dout[31:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:731:26  */
  assign n13569 = mem_dout[32]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:735:26  */
  assign n13570 = stat_mem_rd & valid_mem_rd;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:657:5  */
  always @(posedge clk_i or posedge n13460)
    if (n13460)
      n13571 <= 16'b0000000000000000;
    else
      n13571 <= n13480;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:652:3  */
  assign n13573 = ~n13460;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:657:5  */
  assign n13574 = n13573 ? n13727 : valid_mem_rd;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:657:5  */
  always @(posedge clk_i)
    n13575 <= n13574;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:643:5  */
  always @(posedge clk_i or posedge n13450)
    if (n13450)
      n13582 <= 22'b0000000000000000000000;
    else
      n13582 <= acc_tag;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:643:5  */
  always @(posedge clk_i or posedge n13450)
    if (n13450)
      n13583 <= 4'b0000;
    else
      n13583 <= acc_idx;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:640:5  */
  assign n13584 = {15'b000000000000000, swe_i, n13565, n13560, n13555, n13550};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:640:5  */
  assign n13585 = {tag_mem_rd, acc_idx_ff, 6'b000000};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:684:29  */
  reg [21:0] tag_mem[15:0] ; // memory
  always @(posedge clk_i)
    if (1'b1)
      n13587 <= tag_mem[acc_idx];
  always @(posedge clk_i)
    if (new_i)
      tag_mem[acc_idx] <= acc_tag;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:684:29  */
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:682:17  */
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13589 = acc_idx[3]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13590 = ~n13589;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13591 = acc_idx[2]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13592 = ~n13591;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13593 = n13590 & n13592;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13594 = n13590 & n13591;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13595 = n13589 & n13592;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13596 = n13589 & n13591;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13597 = acc_idx[1]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13598 = ~n13597;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13599 = n13593 & n13598;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13600 = n13593 & n13597;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13601 = n13594 & n13598;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13602 = n13594 & n13597;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13603 = n13595 & n13598;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13604 = n13595 & n13597;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13605 = n13596 & n13598;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13606 = n13596 & n13597;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13607 = acc_idx[0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13608 = ~n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13609 = n13599 & n13608;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13610 = n13599 & n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13611 = n13600 & n13608;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13612 = n13600 & n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13613 = n13601 & n13608;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13614 = n13601 & n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13615 = n13602 & n13608;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13616 = n13602 & n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13617 = n13603 & n13608;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13618 = n13603 & n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13619 = n13604 & n13608;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13620 = n13604 & n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13621 = n13605 & n13608;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13622 = n13605 & n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13623 = n13606 & n13608;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13624 = n13606 & n13607;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:21  */
  assign n13625 = valid_mem[0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13626 = n13609 ? 1'b1 : n13625;
  assign n13627 = valid_mem[1]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13628 = n13610 ? 1'b1 : n13627;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:660:19  */
  assign n13629 = valid_mem[2]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13630 = n13611 ? 1'b1 : n13629;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:652:3  */
  assign n13631 = valid_mem[3]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13632 = n13612 ? 1'b1 : n13631;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:638:3  */
  assign n13633 = valid_mem[4]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13634 = n13613 ? 1'b1 : n13633;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:579:24  */
  assign n13635 = valid_mem[5]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13636 = n13614 ? 1'b1 : n13635;
  assign n13637 = valid_mem[6]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13638 = n13615 ? 1'b1 : n13637;
  assign n13639 = valid_mem[7]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13640 = n13616 ? 1'b1 : n13639;
  assign n13641 = valid_mem[8]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13642 = n13617 ? 1'b1 : n13641;
  assign n13643 = valid_mem[9]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13644 = n13618 ? 1'b1 : n13643;
  assign n13645 = valid_mem[10]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13646 = n13619 ? 1'b1 : n13645;
  assign n13647 = valid_mem[11]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13648 = n13620 ? 1'b1 : n13647;
  assign n13649 = valid_mem[12]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13650 = n13621 ? 1'b1 : n13649;
  assign n13651 = valid_mem[13]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13652 = n13622 ? 1'b1 : n13651;
  assign n13653 = valid_mem[14]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13654 = n13623 ? 1'b1 : n13653;
  assign n13655 = valid_mem[15]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:659:9  */
  assign n13656 = n13624 ? 1'b1 : n13655;
  assign n13657 = {n13656, n13654, n13652, n13650, n13648, n13646, n13644, n13642, n13640, n13638, n13636, n13634, n13632, n13630, n13628, n13626};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13658 = acc_idx[3]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13659 = ~n13658;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13660 = acc_idx[2]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13661 = ~n13660;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13662 = n13659 & n13661;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13663 = n13659 & n13660;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13664 = n13658 & n13661;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13665 = n13658 & n13660;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13666 = acc_idx[1]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13667 = ~n13666;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13668 = n13662 & n13667;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13669 = n13662 & n13666;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13670 = n13663 & n13667;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13671 = n13663 & n13666;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13672 = n13664 & n13667;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13673 = n13664 & n13666;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13674 = n13665 & n13667;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13675 = n13665 & n13666;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13676 = acc_idx[0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13677 = ~n13676;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13678 = n13668 & n13677;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13679 = n13668 & n13676;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13680 = n13669 & n13677;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13681 = n13669 & n13676;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13682 = n13670 & n13677;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13683 = n13670 & n13676;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13684 = n13671 & n13677;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13685 = n13671 & n13676;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13686 = n13672 & n13677;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13687 = n13672 & n13676;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13688 = n13673 & n13677;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13689 = n13673 & n13676;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13690 = n13674 & n13677;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13691 = n13674 & n13676;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13692 = n13675 & n13677;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13693 = n13675 & n13676;
  assign n13694 = valid_mem[0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13695 = n13678 ? 1'b0 : n13694;
  assign n13696 = valid_mem[1]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13697 = n13679 ? 1'b0 : n13696;
  assign n13698 = valid_mem[2]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13699 = n13680 ? 1'b0 : n13698;
  assign n13700 = valid_mem[3]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13701 = n13681 ? 1'b0 : n13700;
  assign n13702 = valid_mem[4]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13703 = n13682 ? 1'b0 : n13702;
  assign n13704 = valid_mem[5]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13705 = n13683 ? 1'b0 : n13704;
  assign n13706 = valid_mem[6]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13707 = n13684 ? 1'b0 : n13706;
  assign n13708 = valid_mem[7]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13709 = n13685 ? 1'b0 : n13708;
  assign n13710 = valid_mem[8]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13711 = n13686 ? 1'b0 : n13710;
  assign n13712 = valid_mem[9]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13713 = n13687 ? 1'b0 : n13712;
  assign n13714 = valid_mem[10]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13715 = n13688 ? 1'b0 : n13714;
  assign n13716 = valid_mem[11]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13717 = n13689 ? 1'b0 : n13716;
  assign n13718 = valid_mem[12]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13719 = n13690 ? 1'b0 : n13718;
  assign n13720 = valid_mem[13]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13721 = n13691 ? 1'b0 : n13720;
  assign n13722 = valid_mem[14]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13723 = n13692 ? 1'b0 : n13722;
  assign n13724 = valid_mem[15]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:663:11  */
  assign n13725 = n13693 ? 1'b0 : n13724;
  assign n13726 = {n13725, n13723, n13721, n13719, n13717, n13715, n13713, n13711, n13709, n13707, n13705, n13703, n13701, n13699, n13697, n13695};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:670:33  */
  assign n13727 = valid_mem[acc_idx * 1 +: 1]; //(Bmux)
endmodule

module neorv32_cache_host_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  rstn_i,
   input  clk_i,
   input  [31:0] \req_i_req_i[addr] ,
   input  [31:0] \req_i_req_i[data] ,
   input  [3:0] \req_i_req_i[ben] ,
   input  \req_i_req_i[stb] ,
   input  \req_i_req_i[rw] ,
   input  \req_i_req_i[src] ,
   input  \req_i_req_i[priv] ,
   input  \req_i_req_i[amo] ,
   input  [3:0] \req_i_req_i[amoop] ,
   input  \req_i_req_i[fence] ,
   input  \req_i_req_i[sleep] ,
   input  \req_i_req_i[debug] ,
   input  bus_busy_i,
   input  hit_i,
   input  [31:0] rdata_i,
   input  rstat_i,
   output [31:0] \rsp_o_rsp_o[data] ,
   output \rsp_o_rsp_o[ack] ,
   output \rsp_o_rsp_o[err] ,
   output bus_sync_o,
   output bus_miss_o,
   output dirty_o,
   output [31:0] addr_o,
   output [3:0] we_o,
   output swe_o,
   output [31:0] wdata_o,
   output wstat_o);
  wire [79:0] n13318;
  wire [31:0] n13320;
  wire n13321;
  wire n13322;
  wire [9:0] ctrl;
  wire n13332;
  wire [2:0] n13337;
  wire n13338;
  wire n13339;
  wire [2:0] n13351;
  wire n13352;
  wire n13353;
  wire n13354;
  wire n13355;
  wire n13356;
  wire n13357;
  wire [31:0] n13358;
  wire [31:0] n13359;
  wire [2:0] n13360;
  wire n13361;
  wire n13363;
  wire n13364;
  wire n13365;
  wire n13366;
  wire n13368;
  wire [2:0] n13371;
  wire [2:0] n13372;
  wire n13375;
  wire [2:0] n13376;
  wire n13378;
  wire n13381;
  wire [1:0] n13384;
  wire [1:0] n13386;
  wire n13389;
  wire [2:0] n13390;
  wire n13392;
  wire n13394;
  wire [2:0] n13396;
  wire n13398;
  wire n13399;
  wire [2:0] n13401;
  wire n13403;
  wire n13407;
  wire [4:0] n13409;
  reg [31:0] n13411;
  wire n13412;
  reg n13414;
  wire n13415;
  reg n13417;
  reg n13422;
  reg n13425;
  reg [2:0] n13427;
  reg n13428;
  reg n13429;
  localparam n13431 = 1'b0;
  localparam [3:0] n13432 = 4'b0000;
  localparam n13433 = 1'b0;
  localparam n13434 = 1'b0;
  reg n13435;
  reg n13436;
  reg [2:0] n13437;
  wire [9:0] n13438;
  wire [33:0] n13439;
  assign \rsp_o_rsp_o[data]  = n13320; //(module output)
  assign \rsp_o_rsp_o[ack]  = n13321; //(module output)
  assign \rsp_o_rsp_o[err]  = n13322; //(module output)
  assign bus_sync_o = n13422; //(module output)
  assign bus_miss_o = n13425; //(module output)
  assign dirty_o = n13431; //(module output)
  assign addr_o = n13358; //(module output)
  assign we_o = n13432; //(module output)
  assign swe_o = n13433; //(module output)
  assign wdata_o = n13359; //(module output)
  assign wstat_o = n13434; //(module output)
  assign n13318 = {\req_i_req_i[debug] , \req_i_req_i[sleep] , \req_i_req_i[fence] , \req_i_req_i[amoop] , \req_i_req_i[amo] , \req_i_req_i[priv] , \req_i_req_i[src] , \req_i_req_i[rw] , \req_i_req_i[stb] , \req_i_req_i[ben] , \req_i_req_i[data] , \req_i_req_i[addr] };
  assign n13320 = n13439[31:0]; // extract
  assign n13321 = n13439[32]; // extract
  assign n13322 = n13439[33]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:419:10  */
  assign ctrl = n13438; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:427:16  */
  assign n13332 = ~rstn_i;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:432:29  */
  assign n13337 = ctrl[5:3]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:433:29  */
  assign n13338 = ctrl[7]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:434:29  */
  assign n13339 = ctrl[9]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:444:31  */
  assign n13351 = ctrl[2:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:445:31  */
  assign n13352 = ctrl[6]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:445:48  */
  assign n13353 = n13318[68]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:445:39  */
  assign n13354 = n13352 | n13353;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:446:31  */
  assign n13355 = ctrl[8]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:446:49  */
  assign n13356 = n13318[77]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:446:40  */
  assign n13357 = n13355 | n13356;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:450:22  */
  assign n13358 = n13318[31:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:453:22  */
  assign n13359 = n13318[63:32]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:15  */
  assign n13360 = ctrl[2:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:468:18  */
  assign n13361 = ctrl[8]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:471:22  */
  assign n13363 = n13318[68]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:471:42  */
  assign n13364 = ctrl[6]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:471:33  */
  assign n13365 = n13363 | n13364;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:472:21  */
  assign n13366 = n13318[69]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:472:31  */
  assign n13368 = 1'b1 & n13366;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:472:11  */
  assign n13371 = n13368 ? 3'b100 : 3'b001;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:471:9  */
  assign n13372 = n13365 ? n13371 : n13351;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:468:9  */
  assign n13375 = n13361 ? 1'b1 : 1'b0;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:468:9  */
  assign n13376 = n13361 ? 3'b011 : n13372;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:466:7  */
  assign n13378 = n13360 == 3'b000;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:488:29  */
  assign n13381 = ~rstat_i;
  assign n13384 = {rstat_i, n13381};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:483:9  */
  assign n13386 = hit_i ? n13384 : 2'b00;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:483:9  */
  assign n13389 = hit_i ? 1'b0 : 1'b1;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:483:9  */
  assign n13390 = hit_i ? 3'b000 : 3'b010;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:479:7  */
  assign n13392 = n13360 == 3'b001;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:499:24  */
  assign n13394 = ~bus_busy_i;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:499:9  */
  assign n13396 = n13394 ? 3'b000 : n13351;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:496:7  */
  assign n13398 = n13360 == 3'b011;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:505:24  */
  assign n13399 = ~bus_busy_i;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:505:9  */
  assign n13401 = n13399 ? 3'b001 : n13351;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:503:7  */
  assign n13403 = n13360 == 3'b010;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:509:7  */
  assign n13407 = n13360 == 3'b100;
  assign n13409 = {n13407, n13403, n13398, n13392, n13378};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:5  */
  always @*
    case (n13409)
      5'b10000: n13411 = 32'b00000000000000000000000000000000;
      5'b01000: n13411 = 32'b00000000000000000000000000000000;
      5'b00100: n13411 = 32'b00000000000000000000000000000000;
      5'b00010: n13411 = rdata_i;
      5'b00001: n13411 = 32'b00000000000000000000000000000000;
      default: n13411 = 32'b00000000000000000000000000000000;
    endcase
  assign n13412 = n13386[0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:5  */
  always @*
    case (n13409)
      5'b10000: n13414 = 1'b0;
      5'b01000: n13414 = 1'b0;
      5'b00100: n13414 = 1'b0;
      5'b00010: n13414 = n13412;
      5'b00001: n13414 = 1'b0;
      default: n13414 = 1'b0;
    endcase
  assign n13415 = n13386[1]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:5  */
  always @*
    case (n13409)
      5'b10000: n13417 = 1'b1;
      5'b01000: n13417 = 1'b0;
      5'b00100: n13417 = 1'b0;
      5'b00010: n13417 = n13415;
      5'b00001: n13417 = 1'b0;
      default: n13417 = 1'b0;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:5  */
  always @*
    case (n13409)
      5'b10000: n13422 = 1'b0;
      5'b01000: n13422 = 1'b0;
      5'b00100: n13422 = 1'b0;
      5'b00010: n13422 = 1'b0;
      5'b00001: n13422 = n13375;
      default: n13422 = 1'b0;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:5  */
  always @*
    case (n13409)
      5'b10000: n13425 = 1'b0;
      5'b01000: n13425 = 1'b0;
      5'b00100: n13425 = 1'b0;
      5'b00010: n13425 = n13389;
      5'b00001: n13425 = 1'b0;
      default: n13425 = 1'b0;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:5  */
  always @*
    case (n13409)
      5'b10000: n13427 = 3'b000;
      5'b01000: n13427 = n13401;
      5'b00100: n13427 = n13396;
      5'b00010: n13427 = n13390;
      5'b00001: n13427 = n13376;
      default: n13427 = 3'b000;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:5  */
  always @*
    case (n13409)
      5'b10000: n13428 = n13354;
      5'b01000: n13428 = n13354;
      5'b00100: n13428 = n13354;
      5'b00010: n13428 = 1'b0;
      5'b00001: n13428 = n13354;
      default: n13428 = n13354;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:464:5  */
  always @*
    case (n13409)
      5'b10000: n13429 = n13357;
      5'b01000: n13429 = n13357;
      5'b00100: n13429 = 1'b0;
      5'b00010: n13429 = n13357;
      5'b00001: n13429 = n13357;
      default: n13429 = n13357;
    endcase
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:431:5  */
  always @(posedge clk_i or posedge n13332)
    if (n13332)
      n13435 <= 1'b0;
    else
      n13435 <= n13339;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:431:5  */
  always @(posedge clk_i or posedge n13332)
    if (n13332)
      n13436 <= 1'b0;
    else
      n13436 <= n13338;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:431:5  */
  always @(posedge clk_i or posedge n13332)
    if (n13332)
      n13437 <= 3'b000;
    else
      n13437 <= n13337;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:427:5  */
  assign n13438 = {n13429, n13435, n13428, n13436, n13427, n13437};
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:427:5  */
  assign n13439 = {n13417, n13414, n13411};
endmodule

module neorv32_xip_phy
  (input  rstn_i,
   input  clk_i,
   input  spi_clk_en_i,
   input  cf_enable_i,
   input  cf_cpha_i,
   input  cf_cpol_i,
   input  op_start_i,
   input  op_final_i,
   input  op_csen_i,
   input  [3:0] op_nbytes_i,
   input  [71:0] op_wdata_i,
   input  spi_dat_i,
   output op_busy_o,
   output [31:0] op_rdata_o,
   output spi_csn_o,
   output spi_clk_o,
   output spi_dat_o);
  wire [83:0] ctrl;
  wire n13165;
  wire n13172;
  wire [2:0] n13178;
  wire [6:0] n13180;
  wire [2:0] n13182;
  wire [2:0] n13183;
  wire n13185;
  wire [2:0] n13187;
  wire [2:0] n13188;
  wire n13190;
  wire n13191;
  wire n13192;
  wire [2:0] n13196;
  wire [2:0] n13197;
  wire [2:0] n13198;
  wire n13200;
  wire n13201;
  wire n13202;
  wire n13203;
  wire n13204;
  wire n13206;
  wire [2:0] n13207;
  wire [2:0] n13208;
  wire n13210;
  wire n13211;
  wire n13212;
  wire [6:0] n13213;
  wire [6:0] n13215;
  wire n13217;
  wire [7:0] n13218;
  wire [2:0] n13219;
  wire [2:0] n13220;
  wire [7:0] n13221;
  wire [7:0] n13222;
  wire n13224;
  wire [70:0] n13225;
  wire n13226;
  wire [71:0] n13227;
  wire n13235;
  wire n13237;
  wire n13239;
  wire n13240;
  wire n13241;
  wire n13242;
  wire n13243;
  wire n13244;
  wire n13245;
  wire n13246;
  wire n13247;
  wire n13248;
  wire n13249;
  wire n13250;
  wire n13251;
  wire n13253;
  wire n13255;
  wire [2:0] n13256;
  wire n13257;
  wire [74:0] n13258;
  wire [74:0] n13259;
  wire [74:0] n13260;
  wire n13262;
  wire [2:0] n13264;
  wire [2:0] n13265;
  wire n13267;
  wire [6:0] n13269;
  reg n13271;
  reg n13272;
  wire [2:0] n13273;
  reg [2:0] n13274;
  wire [71:0] n13275;
  wire [71:0] n13276;
  reg [71:0] n13277;
  wire [6:0] n13278;
  wire [6:0] n13279;
  reg [6:0] n13280;
  wire n13281;
  wire n13282;
  reg n13283;
  wire n13284;
  reg n13285;
  wire n13287;
  wire n13289;
  wire [83:0] n13290;
  wire [83:0] n13291;
  wire [83:0] n13292;
  wire [83:0] n13300;
  wire [2:0] n13304;
  wire n13306;
  wire [2:0] n13307;
  wire n13309;
  wire n13310;
  wire n13311;
  wire n13313;
  wire [31:0] n13314;
  reg [83:0] n13315;
  reg n13316;
  reg n13317;
  assign op_busy_o = n13311; //(module output)
  assign op_rdata_o = n13314; //(module output)
  assign spi_csn_o = n13316; //(module output)
  assign spi_clk_o = n13317; //(module output)
  assign spi_dat_o = n13313; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:453:10  */
  assign ctrl = n13315; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:461:16  */
  assign n13165 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:470:23  */
  assign n13172 = ~cf_enable_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:479:19  */
  assign n13178 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:485:40  */
  assign n13180 = {op_nbytes_i, 3'b000};
  assign n13182 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:487:13  */
  assign n13183 = op_start_i ? 3'b010 : n13182;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:481:11  */
  assign n13185 = n13178 == 3'b000;
  assign n13187 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:494:13  */
  assign n13188 = spi_clk_en_i ? 3'b011 : n13187;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:491:11  */
  assign n13190 = n13178 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:500:37  */
  assign n13191 = ctrl[83]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:500:28  */
  assign n13192 = ~n13191;
  assign n13196 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:504:13  */
  assign n13197 = op_start_i ? 3'b011 : n13196;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:502:13  */
  assign n13198 = op_final_i ? 3'b000 : n13197;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:498:11  */
  assign n13200 = n13178 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:510:35  */
  assign n13201 = ctrl[83]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:510:26  */
  assign n13202 = ~n13201;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:513:30  */
  assign n13203 = ~cf_cpol_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:511:13  */
  assign n13204 = n13206 ? n13203 : n13317;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:511:13  */
  assign n13206 = cf_cpha_i & spi_clk_en_i;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:720:12  */
  assign n13207 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:511:13  */
  assign n13208 = spi_clk_en_i ? 3'b100 : n13207;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:508:11  */
  assign n13210 = n13178 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:521:46  */
  assign n13211 = cf_cpha_i ^ cf_cpol_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:521:31  */
  assign n13212 = ~n13211;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:523:63  */
  assign n13213 = ctrl[81:75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:523:71  */
  assign n13215 = n13213 - 7'b0000001;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:520:13  */
  assign n13217 = spi_clk_en_i ? n13212 : n13317;
  assign n13218 = {spi_dat_i, n13215};
  assign n13219 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:520:13  */
  assign n13220 = spi_clk_en_i ? 3'b101 : n13219;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:76:3  */
  assign n13221 = ctrl[82:75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:520:13  */
  assign n13222 = spi_clk_en_i ? n13218 : n13221;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:518:11  */
  assign n13224 = n13178 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:530:37  */
  assign n13225 = ctrl[73:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:530:72  */
  assign n13226 = ctrl[82]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:530:65  */
  assign n13227 = {n13225, n13226};
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n13235 = ctrl[81]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n13237 = 1'b0 | n13235;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n13239 = ctrl[80]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n13240 = n13237 | n13239;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n13241 = ctrl[79]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n13242 = n13240 | n13241;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n13243 = ctrl[78]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n13244 = n13242 | n13243;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n13245 = ctrl[77]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n13246 = n13244 | n13245;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n13247 = ctrl[76]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n13248 = n13246 | n13247;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n13249 = ctrl[75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n13250 = n13248 | n13249;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:531:44  */
  assign n13251 = ~n13250;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:535:41  */
  assign n13253 = cf_cpha_i ^ cf_cpol_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:531:15  */
  assign n13255 = n13251 ? cf_cpol_i : n13253;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:531:15  */
  assign n13256 = n13251 ? 3'b110 : 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:529:13  */
  assign n13257 = spi_clk_en_i ? n13255 : n13317;
  assign n13258 = {n13227, n13256};
  assign n13259 = ctrl[74:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:529:13  */
  assign n13260 = spi_clk_en_i ? n13258 : n13259;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:527:11  */
  assign n13262 = n13178 == 3'b101;
  assign n13264 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:542:13  */
  assign n13265 = spi_clk_en_i ? 3'b001 : n13264;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:540:11  */
  assign n13267 = n13178 == 3'b110;
  assign n13269 = {n13267, n13262, n13224, n13210, n13200, n13190, n13185};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:479:9  */
  always @*
    case (n13269)
      7'b1000000: n13271 = n13316;
      7'b0100000: n13271 = n13316;
      7'b0010000: n13271 = n13316;
      7'b0001000: n13271 = n13202;
      7'b0000100: n13271 = n13192;
      7'b0000010: n13271 = n13316;
      7'b0000001: n13271 = 1'b1;
      default: n13271 = n13316;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:479:9  */
  always @*
    case (n13269)
      7'b1000000: n13272 = n13317;
      7'b0100000: n13272 = n13257;
      7'b0010000: n13272 = n13217;
      7'b0001000: n13272 = n13204;
      7'b0000100: n13272 = n13317;
      7'b0000010: n13272 = n13317;
      7'b0000001: n13272 = cf_cpol_i;
      default: n13272 = n13317;
    endcase
  assign n13273 = n13260[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:479:9  */
  always @*
    case (n13269)
      7'b1000000: n13274 = n13265;
      7'b0100000: n13274 = n13273;
      7'b0010000: n13274 = n13220;
      7'b0001000: n13274 = n13208;
      7'b0000100: n13274 = n13198;
      7'b0000010: n13274 = n13188;
      7'b0000001: n13274 = n13183;
      default: n13274 = 3'b000;
    endcase
  assign n13275 = n13260[74:3]; // extract
  assign n13276 = ctrl[74:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:479:9  */
  always @*
    case (n13269)
      7'b1000000: n13277 = n13276;
      7'b0100000: n13277 = n13275;
      7'b0010000: n13277 = n13276;
      7'b0001000: n13277 = n13276;
      7'b0000100: n13277 = n13276;
      7'b0000010: n13277 = op_wdata_i;
      7'b0000001: n13277 = n13276;
      default: n13277 = n13276;
    endcase
  assign n13278 = n13222[6:0]; // extract
  assign n13279 = ctrl[81:75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:479:9  */
  always @*
    case (n13269)
      7'b1000000: n13280 = n13279;
      7'b0100000: n13280 = n13279;
      7'b0010000: n13280 = n13278;
      7'b0001000: n13280 = n13279;
      7'b0000100: n13280 = 7'b0100000;
      7'b0000010: n13280 = n13279;
      7'b0000001: n13280 = n13180;
      default: n13280 = n13279;
    endcase
  assign n13281 = n13222[7]; // extract
  assign n13282 = ctrl[82]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:479:9  */
  always @*
    case (n13269)
      7'b1000000: n13283 = n13282;
      7'b0100000: n13283 = n13282;
      7'b0010000: n13283 = n13281;
      7'b0001000: n13283 = n13282;
      7'b0000100: n13283 = n13282;
      7'b0000010: n13283 = n13282;
      7'b0000001: n13283 = n13282;
      default: n13283 = n13282;
    endcase
  assign n13284 = ctrl[83]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:479:9  */
  always @*
    case (n13269)
      7'b1000000: n13285 = n13284;
      7'b0100000: n13285 = n13284;
      7'b0010000: n13285 = n13284;
      7'b0001000: n13285 = n13284;
      7'b0000100: n13285 = n13284;
      7'b0000010: n13285 = n13284;
      7'b0000001: n13285 = op_csen_i;
      default: n13285 = n13284;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:470:7  */
  assign n13287 = n13172 ? 1'b1 : n13271;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:470:7  */
  assign n13289 = n13172 ? 1'b0 : n13272;
  assign n13290 = {n13285, n13283, n13280, n13277, n13274};
  assign n13291 = {1'b0, 1'b0, 7'b0000000, 72'b000000000000000000000000000000000000000000000000000000000000000000000000, 3'b000};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:470:7  */
  assign n13292 = n13172 ? n13291 : n13290;
  assign n13300 = {1'b0, 1'b0, 7'b0000000, 72'b000000000000000000000000000000000000000000000000000000000000000000000000, 3'b000};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:556:31  */
  assign n13304 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:556:37  */
  assign n13306 = n13304 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:556:56  */
  assign n13307 = ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:556:62  */
  assign n13309 = n13307 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:556:47  */
  assign n13310 = n13306 | n13309;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:556:20  */
  assign n13311 = n13310 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:559:25  */
  assign n13313 = ctrl[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:562:26  */
  assign n13314 = ctrl[34:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:469:5  */
  always @(posedge clk_i or posedge n13165)
    if (n13165)
      n13315 <= n13300;
    else
      n13315 <= n13292;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:469:5  */
  always @(posedge clk_i or posedge n13165)
    if (n13165)
      n13316 <= 1'b1;
    else
      n13316 <= n13287;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:469:5  */
  always @(posedge clk_i or posedge n13165)
    if (n13165)
      n13317 <= 1'b0;
    else
      n13317 <= n13289;
endmodule

module neorv32_cpu_lsu_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk_i,
   input  rstn_i,
   input  \ctrl_i_ctrl_i[if_fence] ,
   input  \ctrl_i_ctrl_i[rf_wb_en] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs1] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs2] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rd] ,
   input  \ctrl_i_ctrl_i[rf_zero_we] ,
   input  [2:0] \ctrl_i_ctrl_i[alu_op] ,
   input  \ctrl_i_ctrl_i[alu_sub] ,
   input  \ctrl_i_ctrl_i[alu_opa_mux] ,
   input  \ctrl_i_ctrl_i[alu_opb_mux] ,
   input  \ctrl_i_ctrl_i[alu_unsigned] ,
   input  \ctrl_i_ctrl_i[alu_cp_alu] ,
   input  \ctrl_i_ctrl_i[alu_cp_cfu] ,
   input  \ctrl_i_ctrl_i[alu_cp_fpu] ,
   input  \ctrl_i_ctrl_i[lsu_req] ,
   input  \ctrl_i_ctrl_i[lsu_rw] ,
   input  \ctrl_i_ctrl_i[lsu_mo_we] ,
   input  \ctrl_i_ctrl_i[lsu_fence] ,
   input  \ctrl_i_ctrl_i[lsu_priv] ,
   input  [2:0] \ctrl_i_ctrl_i[ir_funct3] ,
   input  [11:0] \ctrl_i_ctrl_i[ir_funct12] ,
   input  [6:0] \ctrl_i_ctrl_i[ir_opcode] ,
   input  \ctrl_i_ctrl_i[cpu_priv] ,
   input  \ctrl_i_ctrl_i[cpu_sleep] ,
   input  \ctrl_i_ctrl_i[cpu_trap] ,
   input  \ctrl_i_ctrl_i[cpu_debug] ,
   input  [31:0] addr_i,
   input  [31:0] wdata_i,
   input  pmp_fault_i,
   input  [31:0] \dbus_rsp_i_dbus_rsp_i[data] ,
   input  \dbus_rsp_i_dbus_rsp_i[ack] ,
   input  \dbus_rsp_i_dbus_rsp_i[err] ,
   output [31:0] rdata_o,
   output [31:0] mar_o,
   output wait_o,
   output [3:0] err_o,
   output [31:0] \dbus_req_o_dbus_req_o[addr] ,
   output [31:0] \dbus_req_o_dbus_req_o[data] ,
   output [3:0] \dbus_req_o_dbus_req_o[ben] ,
   output \dbus_req_o_dbus_req_o[stb] ,
   output \dbus_req_o_dbus_req_o[rw] ,
   output \dbus_req_o_dbus_req_o[src] ,
   output \dbus_req_o_dbus_req_o[priv] ,
   output \dbus_req_o_dbus_req_o[amo] ,
   output [3:0] \dbus_req_o_dbus_req_o[amoop] ,
   output \dbus_req_o_dbus_req_o[fence] ,
   output \dbus_req_o_dbus_req_o[sleep] ,
   output \dbus_req_o_dbus_req_o[debug] );
  wire [58:0] n12804;
  wire [31:0] n12810;
  wire [31:0] n12811;
  wire [3:0] n12812;
  wire n12813;
  wire n12814;
  wire n12815;
  wire n12816;
  wire n12817;
  wire [3:0] n12818;
  wire n12819;
  wire n12820;
  wire n12821;
  wire [33:0] n12822;
  wire [31:0] mar;
  wire misaligned;
  wire arbiter_req;
  wire arbiter_err;
  wire [3:0] amo_cmd;
  wire n12824;
  wire n12826;
  wire [1:0] n12827;
  wire n12829;
  wire n12830;
  wire n12832;
  wire n12833;
  wire n12834;
  wire n12835;
  wire [1:0] n12836;
  reg n12838;
  wire n12849;
  wire n12857;
  wire n12858;
  wire n12859;
  wire n12861;
  wire n12863;
  wire [1:0] n12864;
  wire [7:0] n12865;
  wire [7:0] n12866;
  wire [15:0] n12867;
  wire [7:0] n12868;
  wire [23:0] n12869;
  wire [7:0] n12870;
  wire [31:0] n12871;
  wire n12872;
  wire n12873;
  wire n12874;
  wire n12875;
  wire n12876;
  wire n12877;
  wire n12878;
  wire n12879;
  wire n12880;
  wire n12881;
  wire n12882;
  wire n12883;
  wire n12884;
  wire n12885;
  wire n12886;
  wire n12887;
  wire n12889;
  wire [15:0] n12890;
  wire [15:0] n12891;
  wire [31:0] n12892;
  wire n12893;
  wire n12894;
  wire [1:0] n12895;
  wire n12896;
  wire n12897;
  wire [2:0] n12898;
  wire n12899;
  wire n12900;
  wire [3:0] n12901;
  wire n12903;
  localparam [3:0] n12904 = 4'b1111;
  wire [1:0] n12905;
  reg [31:0] n12906;
  wire n12907;
  wire n12908;
  reg n12909;
  wire n12910;
  wire n12911;
  reg n12912;
  wire n12913;
  wire n12914;
  reg n12915;
  wire n12916;
  wire n12917;
  reg n12918;
  wire [35:0] n12919;
  wire [5:0] n12920;
  wire [35:0] n12933;
  wire [5:0] n12934;
  wire n12940;
  wire n12941;
  wire n12942;
  wire n12947;
  wire [1:0] n12949;
  wire [1:0] n12950;
  wire n12952;
  wire n12953;
  wire n12954;
  wire n12955;
  wire [3:0] n12961;
  wire [3:0] n12962;
  wire [3:0] n12963;
  wire [3:0] n12964;
  wire [3:0] n12965;
  wire [3:0] n12966;
  wire [15:0] n12967;
  wire [7:0] n12968;
  wire [23:0] n12969;
  wire [7:0] n12971;
  wire [31:0] n12972;
  wire n12974;
  wire n12976;
  wire n12977;
  wire n12978;
  wire n12979;
  wire [3:0] n12985;
  wire [3:0] n12986;
  wire [3:0] n12987;
  wire [3:0] n12988;
  wire [3:0] n12989;
  wire [3:0] n12990;
  wire [15:0] n12991;
  wire [7:0] n12992;
  wire [23:0] n12993;
  wire [7:0] n12995;
  wire [31:0] n12996;
  wire n12998;
  wire n13000;
  wire n13001;
  wire n13002;
  wire n13003;
  wire [3:0] n13009;
  wire [3:0] n13010;
  wire [3:0] n13011;
  wire [3:0] n13012;
  wire [3:0] n13013;
  wire [3:0] n13014;
  wire [15:0] n13015;
  wire [7:0] n13016;
  wire [23:0] n13017;
  wire [7:0] n13019;
  wire [31:0] n13020;
  wire n13022;
  wire n13024;
  wire n13025;
  wire n13026;
  wire n13027;
  wire [3:0] n13033;
  wire [3:0] n13034;
  wire [3:0] n13035;
  wire [3:0] n13036;
  wire [3:0] n13037;
  wire [3:0] n13038;
  wire [15:0] n13039;
  wire [7:0] n13040;
  wire [23:0] n13041;
  wire [7:0] n13043;
  wire [31:0] n13044;
  wire [2:0] n13045;
  reg [31:0] n13046;
  wire n13048;
  wire n13049;
  wire n13050;
  wire n13052;
  wire n13053;
  wire n13054;
  wire n13055;
  wire [3:0] n13061;
  wire [3:0] n13062;
  wire [3:0] n13063;
  wire [3:0] n13064;
  wire [15:0] n13065;
  wire [15:0] n13067;
  wire [31:0] n13068;
  wire n13070;
  wire n13071;
  wire n13072;
  wire n13073;
  wire [3:0] n13079;
  wire [3:0] n13080;
  wire [3:0] n13081;
  wire [3:0] n13082;
  wire [15:0] n13083;
  wire [15:0] n13085;
  wire [31:0] n13086;
  wire [31:0] n13087;
  wire n13089;
  wire [31:0] n13090;
  wire [1:0] n13091;
  reg [31:0] n13092;
  wire [31:0] n13094;
  wire n13101;
  wire n13103;
  wire n13104;
  wire n13105;
  wire n13106;
  wire n13107;
  wire n13108;
  wire n13109;
  wire n13111;
  wire n13112;
  wire n13120;
  wire n13121;
  wire n13122;
  wire n13123;
  wire n13124;
  wire n13125;
  wire n13126;
  wire n13127;
  wire n13128;
  wire n13129;
  wire n13130;
  wire n13131;
  wire n13132;
  wire n13133;
  wire n13134;
  wire n13135;
  wire n13136;
  wire n13137;
  wire n13138;
  wire n13139;
  wire n13140;
  wire [31:0] n13141;
  reg [31:0] n13142;
  wire n13143;
  reg n13144;
  reg n13145;
  reg n13146;
  reg [31:0] n13147;
  wire [3:0] n13148;
  wire [5:0] n13149;
  wire [5:0] n13150;
  reg [5:0] n13151;
  wire n13152;
  wire n13153;
  reg n13154;
  wire [35:0] n13155;
  wire [35:0] n13156;
  reg [35:0] n13157;
  wire [79:0] n13158;
  assign rdata_o = n13147; //(module output)
  assign mar_o = mar; //(module output)
  assign wait_o = n13121; //(module output)
  assign err_o = n13148; //(module output)
  assign \dbus_req_o_dbus_req_o[addr]  = n12810; //(module output)
  assign \dbus_req_o_dbus_req_o[data]  = n12811; //(module output)
  assign \dbus_req_o_dbus_req_o[ben]  = n12812; //(module output)
  assign \dbus_req_o_dbus_req_o[stb]  = n12813; //(module output)
  assign \dbus_req_o_dbus_req_o[rw]  = n12814; //(module output)
  assign \dbus_req_o_dbus_req_o[src]  = n12815; //(module output)
  assign \dbus_req_o_dbus_req_o[priv]  = n12816; //(module output)
  assign \dbus_req_o_dbus_req_o[amo]  = n12817; //(module output)
  assign \dbus_req_o_dbus_req_o[amoop]  = n12818; //(module output)
  assign \dbus_req_o_dbus_req_o[fence]  = n12819; //(module output)
  assign \dbus_req_o_dbus_req_o[sleep]  = n12820; //(module output)
  assign \dbus_req_o_dbus_req_o[debug]  = n12821; //(module output)
  assign n12804 = {\ctrl_i_ctrl_i[cpu_debug] , \ctrl_i_ctrl_i[cpu_trap] , \ctrl_i_ctrl_i[cpu_sleep] , \ctrl_i_ctrl_i[cpu_priv] , \ctrl_i_ctrl_i[ir_opcode] , \ctrl_i_ctrl_i[ir_funct12] , \ctrl_i_ctrl_i[ir_funct3] , \ctrl_i_ctrl_i[lsu_priv] , \ctrl_i_ctrl_i[lsu_fence] , \ctrl_i_ctrl_i[lsu_mo_we] , \ctrl_i_ctrl_i[lsu_rw] , \ctrl_i_ctrl_i[lsu_req] , \ctrl_i_ctrl_i[alu_cp_fpu] , \ctrl_i_ctrl_i[alu_cp_cfu] , \ctrl_i_ctrl_i[alu_cp_alu] , \ctrl_i_ctrl_i[alu_unsigned] , \ctrl_i_ctrl_i[alu_opb_mux] , \ctrl_i_ctrl_i[alu_opa_mux] , \ctrl_i_ctrl_i[alu_sub] , \ctrl_i_ctrl_i[alu_op] , \ctrl_i_ctrl_i[rf_zero_we] , \ctrl_i_ctrl_i[rf_rd] , \ctrl_i_ctrl_i[rf_rs2] , \ctrl_i_ctrl_i[rf_rs1] , \ctrl_i_ctrl_i[rf_wb_en] , \ctrl_i_ctrl_i[if_fence] };
  assign n12810 = n13158[31:0]; // extract
  assign n12811 = n13158[63:32]; // extract
  assign n12812 = n13158[67:64]; // extract
  assign n12813 = n13158[68]; // extract
  assign n12814 = n13158[69]; // extract
  assign n12815 = n13158[70]; // extract
  assign n12816 = n13158[71]; // extract
  assign n12817 = n13158[72]; // extract
  assign n12818 = n13158[76:73]; // extract
  assign n12819 = n13158[77]; // extract
  assign n12820 = n13158[78]; // extract
  assign n12821 = n13158[79]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1026:14  */
  assign n12822 = {\dbus_rsp_i_dbus_rsp_i[err] , \dbus_rsp_i_dbus_rsp_i[ack] , \dbus_rsp_i_dbus_rsp_i[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:42:10  */
  assign mar = n13142; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:43:10  */
  assign misaligned = n13144; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:44:10  */
  assign arbiter_req = n13145; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:45:10  */
  assign arbiter_err = n13146; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:46:10  */
  assign amo_cmd = 4'b0000; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:54:16  */
  assign n12824 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:58:18  */
  assign n12826 = n12804[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:60:30  */
  assign n12827 = n12804[34:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:61:11  */
  assign n12829 = n12827 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:62:46  */
  assign n12830 = addr_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:62:11  */
  assign n12832 = n12827 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:63:46  */
  assign n12833 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:63:59  */
  assign n12834 = addr_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:63:50  */
  assign n12835 = n12833 | n12834;
  assign n12836 = {n12832, n12829};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:60:9  */
  always @*
    case (n12836)
      2'b10: n12838 = n12830;
      2'b01: n12838 = 1'b0;
      default: n12838 = n12835;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:78:16  */
  assign n12849 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:86:18  */
  assign n12857 = n12804[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:88:36  */
  assign n12858 = n12804[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:89:36  */
  assign n12859 = n12804[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:90:74  */
  assign n12861 = n12804[50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:90:54  */
  assign n12863 = 1'b0 & n12861;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:93:30  */
  assign n12864 = n12804[34:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:95:41  */
  assign n12865 = wdata_i[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:95:63  */
  assign n12866 = wdata_i[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:95:54  */
  assign n12867 = {n12865, n12866};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:95:85  */
  assign n12868 = wdata_i[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:95:76  */
  assign n12869 = {n12867, n12868};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:95:107  */
  assign n12870 = wdata_i[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:95:98  */
  assign n12871 = {n12869, n12870};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:96:45  */
  assign n12872 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:96:35  */
  assign n12873 = ~n12872;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:96:65  */
  assign n12874 = addr_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:96:55  */
  assign n12875 = ~n12874;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:96:50  */
  assign n12876 = n12873 & n12875;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:97:45  */
  assign n12877 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:97:35  */
  assign n12878 = ~n12877;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:97:65  */
  assign n12879 = addr_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:97:50  */
  assign n12880 = n12878 & n12879;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:98:45  */
  assign n12881 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:98:65  */
  assign n12882 = addr_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:98:55  */
  assign n12883 = ~n12882;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:98:50  */
  assign n12884 = n12881 & n12883;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:99:45  */
  assign n12885 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:99:65  */
  assign n12886 = addr_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:99:50  */
  assign n12887 = n12885 & n12886;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:94:11  */
  assign n12889 = n12864 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:101:39  */
  assign n12890 = wdata_i[15:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:101:62  */
  assign n12891 = wdata_i[15:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:101:53  */
  assign n12892 = {n12890, n12891};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:38  */
  assign n12893 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:50  */
  assign n12894 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:42  */
  assign n12895 = {n12893, n12894};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:67  */
  assign n12896 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:57  */
  assign n12897 = ~n12896;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:54  */
  assign n12898 = {n12895, n12897};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:85  */
  assign n12899 = addr_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:75  */
  assign n12900 = ~n12899;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:102:72  */
  assign n12901 = {n12898, n12900};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:100:11  */
  assign n12903 = n12864 == 2'b01;
  assign n12905 = {n12903, n12889};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:93:9  */
  always @*
    case (n12905)
      2'b10: n12906 = n12892;
      2'b01: n12906 = n12871;
      default: n12906 = wdata_i;
    endcase
  assign n12907 = n12901[0]; // extract
  assign n12908 = n12904[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:93:9  */
  always @*
    case (n12905)
      2'b10: n12909 = n12907;
      2'b01: n12909 = n12876;
      default: n12909 = n12908;
    endcase
  assign n12910 = n12901[1]; // extract
  assign n12911 = n12904[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:93:9  */
  always @*
    case (n12905)
      2'b10: n12912 = n12910;
      2'b01: n12912 = n12880;
      default: n12912 = n12911;
    endcase
  assign n12913 = n12901[2]; // extract
  assign n12914 = n12904[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:93:9  */
  always @*
    case (n12905)
      2'b10: n12915 = n12913;
      2'b01: n12915 = n12884;
      default: n12915 = n12914;
    endcase
  assign n12916 = n12901[3]; // extract
  assign n12917 = n12904[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:93:9  */
  always @*
    case (n12905)
      2'b10: n12918 = n12916;
      2'b01: n12918 = n12887;
      default: n12918 = n12917;
    endcase
  assign n12919 = {n12918, n12915, n12912, n12909, n12906};
  assign n12920 = {amo_cmd, n12863, n12859};
  assign n12933 = {4'b0000, 32'b00000000000000000000000000000000};
  assign n12934 = {4'b0000, 1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:112:30  */
  assign n12940 = n12804[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:113:30  */
  assign n12941 = n12804[56]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:114:30  */
  assign n12942 = n12804[58]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:141:16  */
  assign n12947 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:146:30  */
  assign n12949 = n12804[34:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:148:21  */
  assign n12950 = mar[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:149:74  */
  assign n12952 = n12804[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:149:54  */
  assign n12953 = ~n12952;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:149:98  */
  assign n12954 = n12822[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:149:79  */
  assign n12955 = n12953 & n12954;
  assign n12961 = {n12955, n12955, n12955, n12955};
  assign n12962 = {n12955, n12955, n12955, n12955};
  assign n12963 = {n12955, n12955, n12955, n12955};
  assign n12964 = {n12955, n12955, n12955, n12955};
  assign n12965 = {n12955, n12955, n12955, n12955};
  assign n12966 = {n12955, n12955, n12955, n12955};
  assign n12967 = {n12961, n12962, n12963, n12964};
  assign n12968 = {n12965, n12966};
  assign n12969 = {n12967, n12968};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:149:125  */
  assign n12971 = n12822[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:149:108  */
  assign n12972 = {n12969, n12971};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:149:15  */
  assign n12974 = n12950 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:150:74  */
  assign n12976 = n12804[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:150:54  */
  assign n12977 = ~n12976;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:150:98  */
  assign n12978 = n12822[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:150:79  */
  assign n12979 = n12977 & n12978;
  assign n12985 = {n12979, n12979, n12979, n12979};
  assign n12986 = {n12979, n12979, n12979, n12979};
  assign n12987 = {n12979, n12979, n12979, n12979};
  assign n12988 = {n12979, n12979, n12979, n12979};
  assign n12989 = {n12979, n12979, n12979, n12979};
  assign n12990 = {n12979, n12979, n12979, n12979};
  assign n12991 = {n12985, n12986, n12987, n12988};
  assign n12992 = {n12989, n12990};
  assign n12993 = {n12991, n12992};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:150:125  */
  assign n12995 = n12822[15:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:150:108  */
  assign n12996 = {n12993, n12995};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:150:15  */
  assign n12998 = n12950 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:151:74  */
  assign n13000 = n12804[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:151:54  */
  assign n13001 = ~n13000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:151:98  */
  assign n13002 = n12822[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:151:79  */
  assign n13003 = n13001 & n13002;
  assign n13009 = {n13003, n13003, n13003, n13003};
  assign n13010 = {n13003, n13003, n13003, n13003};
  assign n13011 = {n13003, n13003, n13003, n13003};
  assign n13012 = {n13003, n13003, n13003, n13003};
  assign n13013 = {n13003, n13003, n13003, n13003};
  assign n13014 = {n13003, n13003, n13003, n13003};
  assign n13015 = {n13009, n13010, n13011, n13012};
  assign n13016 = {n13013, n13014};
  assign n13017 = {n13015, n13016};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:151:125  */
  assign n13019 = n12822[23:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:151:108  */
  assign n13020 = {n13017, n13019};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:151:15  */
  assign n13022 = n12950 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:152:74  */
  assign n13024 = n12804[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:152:54  */
  assign n13025 = ~n13024;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:152:98  */
  assign n13026 = n12822[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:152:79  */
  assign n13027 = n13025 & n13026;
  assign n13033 = {n13027, n13027, n13027, n13027};
  assign n13034 = {n13027, n13027, n13027, n13027};
  assign n13035 = {n13027, n13027, n13027, n13027};
  assign n13036 = {n13027, n13027, n13027, n13027};
  assign n13037 = {n13027, n13027, n13027, n13027};
  assign n13038 = {n13027, n13027, n13027, n13027};
  assign n13039 = {n13033, n13034, n13035, n13036};
  assign n13040 = {n13037, n13038};
  assign n13041 = {n13039, n13040};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:152:125  */
  assign n13043 = n12822[31:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:152:108  */
  assign n13044 = {n13041, n13043};
  assign n13045 = {n13022, n12998, n12974};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:148:13  */
  always @*
    case (n13045)
      3'b100: n13046 = n13020;
      3'b010: n13046 = n12996;
      3'b001: n13046 = n12972;
      default: n13046 = n13044;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:147:11  */
  assign n13048 = n12949 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:155:20  */
  assign n13049 = mar[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:155:24  */
  assign n13050 = ~n13049;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:156:59  */
  assign n13052 = n12804[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:156:39  */
  assign n13053 = ~n13052;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:156:83  */
  assign n13054 = n12822[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:156:64  */
  assign n13055 = n13053 & n13054;
  assign n13061 = {n13055, n13055, n13055, n13055};
  assign n13062 = {n13055, n13055, n13055, n13055};
  assign n13063 = {n13055, n13055, n13055, n13055};
  assign n13064 = {n13055, n13055, n13055, n13055};
  assign n13065 = {n13061, n13062, n13063, n13064};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:156:110  */
  assign n13067 = n12822[15:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:156:93  */
  assign n13068 = {n13065, n13067};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:158:59  */
  assign n13070 = n12804[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:158:39  */
  assign n13071 = ~n13070;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:158:83  */
  assign n13072 = n12822[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:158:64  */
  assign n13073 = n13071 & n13072;
  assign n13079 = {n13073, n13073, n13073, n13073};
  assign n13080 = {n13073, n13073, n13073, n13073};
  assign n13081 = {n13073, n13073, n13073, n13073};
  assign n13082 = {n13073, n13073, n13073, n13073};
  assign n13083 = {n13079, n13080, n13081, n13082};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:158:110  */
  assign n13085 = n12822[31:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:158:93  */
  assign n13086 = {n13083, n13085};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:155:13  */
  assign n13087 = n13050 ? n13068 : n13086;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:154:11  */
  assign n13089 = n12949 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:161:35  */
  assign n13090 = n12822[31:0]; // extract
  assign n13091 = {n13089, n13048};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:146:9  */
  always @*
    case (n13091)
      2'b10: n13092 = n13087;
      2'b01: n13092 = n13046;
      default: n13092 = n13090;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:145:7  */
  assign n13094 = arbiter_req ? n13092 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:172:16  */
  assign n13101 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:176:33  */
  assign n13103 = n12822[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:176:37  */
  assign n13104 = n13103 | pmp_fault_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:177:23  */
  assign n13105 = ~arbiter_req;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:178:31  */
  assign n13106 = n12804[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:179:25  */
  assign n13107 = n12822[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:179:47  */
  assign n13108 = n12804[57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:179:36  */
  assign n13109 = n13107 | n13108;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:179:7  */
  assign n13111 = n13109 ? 1'b0 : arbiter_req;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:177:7  */
  assign n13112 = n13105 ? n13106 : n13111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:186:28  */
  assign n13120 = n12822[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:186:13  */
  assign n13121 = ~n13120;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:189:43  */
  assign n13122 = n12804[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:189:32  */
  assign n13123 = ~n13122;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:189:27  */
  assign n13124 = arbiter_req & n13123;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:189:51  */
  assign n13125 = n13124 & misaligned;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:190:43  */
  assign n13126 = n12804[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:190:32  */
  assign n13127 = ~n13126;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:190:27  */
  assign n13128 = arbiter_req & n13127;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:190:51  */
  assign n13129 = n13128 & arbiter_err;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:191:43  */
  assign n13130 = n12804[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:191:27  */
  assign n13131 = arbiter_req & n13130;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:191:51  */
  assign n13132 = n13131 & misaligned;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:192:43  */
  assign n13133 = n12804[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:192:27  */
  assign n13134 = arbiter_req & n13133;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:192:51  */
  assign n13135 = n13134 & arbiter_err;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:195:28  */
  assign n13136 = n12804[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:195:41  */
  assign n13137 = ~misaligned;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:195:36  */
  assign n13138 = n13136 & n13137;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:195:62  */
  assign n13139 = ~pmp_fault_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:195:57  */
  assign n13140 = n13138 & n13139;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:57:5  */
  assign n13141 = n12826 ? addr_i : mar;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:57:5  */
  always @(posedge clk_i or posedge n12824)
    if (n12824)
      n13142 <= 32'b00000000000000000000000000000000;
    else
      n13142 <= n13141;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:57:5  */
  assign n13143 = n12826 ? n12838 : misaligned;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:57:5  */
  always @(posedge clk_i or posedge n12824)
    if (n12824)
      n13144 <= 1'b0;
    else
      n13144 <= n13143;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:175:5  */
  always @(posedge clk_i or posedge n13101)
    if (n13101)
      n13145 <= 1'b0;
    else
      n13145 <= n13112;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:175:5  */
  always @(posedge clk_i or posedge n13101)
    if (n13101)
      n13146 <= 1'b0;
    else
      n13146 <= n13104;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:143:5  */
  always @(posedge clk_i or posedge n12947)
    if (n12947)
      n13147 <= 32'b00000000000000000000000000000000;
    else
      n13147 <= n13094;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:141:5  */
  assign n13148 = {n13135, n13132, n13129, n13125};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  assign n13149 = n13158[76:71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  assign n13150 = n12857 ? n12920 : n13149;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  always @(posedge clk_i or posedge n12849)
    if (n12849)
      n13151 <= n12934;
    else
      n13151 <= n13150;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  assign n13152 = n13158[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  assign n13153 = n12857 ? n12858 : n13152;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  always @(posedge clk_i or posedge n12849)
    if (n12849)
      n13154 <= 1'b0;
    else
      n13154 <= n13153;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  assign n13155 = n13158[67:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  assign n13156 = n12857 ? n12919 : n13155;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:85:5  */
  always @(posedge clk_i or posedge n12849)
    if (n12849)
      n13157 <= n12933;
    else
      n13157 <= n13156;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_lsu.vhd:78:5  */
  assign n13158 = {n12942, n12941, n12940, n13151, 1'b0, n13154, n13140, n13157, mar};
endmodule

module neorv32_cpu_alu_f8bf199495d218f30da53ac11031539acc71c5ae
  (input  clk_i,
   input  rstn_i,
   input  \ctrl_i_ctrl_i[if_fence] ,
   input  \ctrl_i_ctrl_i[rf_wb_en] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs1] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs2] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rd] ,
   input  \ctrl_i_ctrl_i[rf_zero_we] ,
   input  [2:0] \ctrl_i_ctrl_i[alu_op] ,
   input  \ctrl_i_ctrl_i[alu_sub] ,
   input  \ctrl_i_ctrl_i[alu_opa_mux] ,
   input  \ctrl_i_ctrl_i[alu_opb_mux] ,
   input  \ctrl_i_ctrl_i[alu_unsigned] ,
   input  \ctrl_i_ctrl_i[alu_cp_alu] ,
   input  \ctrl_i_ctrl_i[alu_cp_cfu] ,
   input  \ctrl_i_ctrl_i[alu_cp_fpu] ,
   input  \ctrl_i_ctrl_i[lsu_req] ,
   input  \ctrl_i_ctrl_i[lsu_rw] ,
   input  \ctrl_i_ctrl_i[lsu_mo_we] ,
   input  \ctrl_i_ctrl_i[lsu_fence] ,
   input  \ctrl_i_ctrl_i[lsu_priv] ,
   input  [2:0] \ctrl_i_ctrl_i[ir_funct3] ,
   input  [11:0] \ctrl_i_ctrl_i[ir_funct12] ,
   input  [6:0] \ctrl_i_ctrl_i[ir_opcode] ,
   input  \ctrl_i_ctrl_i[cpu_priv] ,
   input  \ctrl_i_ctrl_i[cpu_sleep] ,
   input  \ctrl_i_ctrl_i[cpu_trap] ,
   input  \ctrl_i_ctrl_i[cpu_debug] ,
   input  csr_we_i,
   input  [11:0] csr_addr_i,
   input  [31:0] csr_wdata_i,
   input  [31:0] rs1_i,
   input  [31:0] rs2_i,
   input  [31:0] rs3_i,
   input  [31:0] pc_i,
   input  [31:0] imm_i,
   output [31:0] csr_rdata_o,
   output [1:0] cmp_o,
   output [31:0] res_o,
   output [31:0] add_o,
   output cp_done_o);
  wire [58:0] n12604;
  wire [32:0] cmp_rs1;
  wire [32:0] cmp_rs2;
  wire [1:0] cmp;
  wire [31:0] opa;
  wire [31:0] opb;
  wire [32:0] opa_x;
  wire [32:0] opb_x;
  wire [32:0] addsub_res;
  wire [31:0] cp_res;
  wire [223:0] cp_result;
  wire [6:0] cp_valid;
  wire [4:0] cp_shamt;
  wire [31:0] csr_rdata_fpu;
  wire [31:0] csr_rdata_cfu;
  wire n12610;
  wire n12611;
  wire n12612;
  wire n12613;
  wire [32:0] n12614;
  wire n12615;
  wire n12616;
  wire n12617;
  wire n12618;
  wire [32:0] n12619;
  wire n12621;
  wire n12622;
  wire n12625;
  wire n12626;
  wire n12628;
  wire [31:0] n12629;
  wire n12630;
  wire [31:0] n12631;
  wire n12632;
  wire n12633;
  wire n12634;
  wire n12635;
  wire [32:0] n12636;
  wire n12637;
  wire n12638;
  wire n12639;
  wire n12640;
  wire [32:0] n12641;
  wire [32:0] n12642;
  wire n12643;
  wire [32:0] n12644;
  wire [32:0] n12645;
  wire [31:0] n12646;
  wire [2:0] n12648;
  wire n12650;
  wire [31:0] n12651;
  wire n12653;
  wire n12655;
  wire n12656;
  wire n12658;
  wire n12660;
  wire [31:0] n12661;
  wire n12663;
  wire [31:0] n12664;
  wire n12666;
  wire [31:0] n12667;
  wire n12669;
  wire [7:0] n12670;
  wire n12672;
  wire n12673;
  wire n12674;
  wire n12675;
  wire n12676;
  wire n12677;
  reg n12679;
  wire [30:0] n12681;
  wire [30:0] n12682;
  wire [30:0] n12683;
  wire [30:0] n12684;
  wire [30:0] n12685;
  wire [30:0] n12686;
  reg [30:0] n12689;
  wire n12693;
  wire n12694;
  wire n12695;
  wire n12696;
  wire n12697;
  wire n12698;
  wire n12699;
  wire n12700;
  wire n12701;
  wire n12702;
  wire n12703;
  wire n12704;
  wire n12705;
  wire [31:0] n12706;
  wire [31:0] n12707;
  wire [31:0] n12708;
  wire [31:0] n12709;
  wire [31:0] n12710;
  wire [31:0] n12711;
  wire [31:0] n12712;
  wire [31:0] n12713;
  wire [31:0] n12714;
  wire [31:0] n12715;
  wire [31:0] n12716;
  wire [31:0] n12717;
  wire [31:0] n12718;
  wire [31:0] n12719;
  wire [4:0] n12721;
  wire [31:0] \neorv32_cpu_cp_shifter_inst.res_o ;
  wire \neorv32_cpu_cp_shifter_inst.valid_o ;
  wire n12722;
  wire n12723;
  wire [4:0] n12724;
  wire [4:0] n12725;
  wire [4:0] n12726;
  wire n12727;
  wire [2:0] n12728;
  wire n12729;
  wire n12730;
  wire n12731;
  wire n12732;
  wire n12733;
  wire n12734;
  wire n12735;
  wire n12736;
  wire n12737;
  wire n12738;
  wire n12739;
  wire n12740;
  wire [2:0] n12741;
  wire [11:0] n12742;
  wire [6:0] n12743;
  wire n12744;
  wire n12745;
  wire n12746;
  wire n12747;
  wire [31:0] \neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst.res_o ;
  wire \neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst.valid_o ;
  wire n12750;
  wire n12751;
  wire [4:0] n12752;
  wire [4:0] n12753;
  wire [4:0] n12754;
  wire n12755;
  wire [2:0] n12756;
  wire n12757;
  wire n12758;
  wire n12759;
  wire n12760;
  wire n12761;
  wire n12762;
  wire n12763;
  wire n12764;
  wire n12765;
  wire n12766;
  wire n12767;
  wire n12768;
  wire [2:0] n12769;
  wire [11:0] n12770;
  wire [6:0] n12771;
  wire n12772;
  wire n12773;
  wire n12774;
  wire n12775;
  wire [1:0] n12796;
  wire [223:0] n12797;
  wire [6:0] n12798;
  wire [31:0] n12803;
  assign csr_rdata_o = n12719; //(module output)
  assign cmp_o = cmp; //(module output)
  assign res_o = n12803; //(module output)
  assign add_o = n12646; //(module output)
  assign cp_done_o = n12705; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:130:27  */
  assign n12604 = {\ctrl_i_ctrl_i[cpu_debug] , \ctrl_i_ctrl_i[cpu_trap] , \ctrl_i_ctrl_i[cpu_sleep] , \ctrl_i_ctrl_i[cpu_priv] , \ctrl_i_ctrl_i[ir_opcode] , \ctrl_i_ctrl_i[ir_funct12] , \ctrl_i_ctrl_i[ir_funct3] , \ctrl_i_ctrl_i[lsu_priv] , \ctrl_i_ctrl_i[lsu_fence] , \ctrl_i_ctrl_i[lsu_mo_we] , \ctrl_i_ctrl_i[lsu_rw] , \ctrl_i_ctrl_i[lsu_req] , \ctrl_i_ctrl_i[alu_cp_fpu] , \ctrl_i_ctrl_i[alu_cp_cfu] , \ctrl_i_ctrl_i[alu_cp_alu] , \ctrl_i_ctrl_i[alu_unsigned] , \ctrl_i_ctrl_i[alu_opb_mux] , \ctrl_i_ctrl_i[alu_opa_mux] , \ctrl_i_ctrl_i[alu_sub] , \ctrl_i_ctrl_i[alu_op] , \ctrl_i_ctrl_i[rf_zero_we] , \ctrl_i_ctrl_i[rf_rd] , \ctrl_i_ctrl_i[rf_rs2] , \ctrl_i_ctrl_i[rf_rs1] , \ctrl_i_ctrl_i[rf_wb_en] , \ctrl_i_ctrl_i[if_fence] };
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:69:10  */
  assign cmp_rs1 = n12614; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:70:10  */
  assign cmp_rs2 = n12619; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:71:10  */
  assign cmp = n12796; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:74:10  */
  assign opa = n12629; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:74:17  */
  assign opb = n12631; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:75:10  */
  assign opa_x = n12636; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:75:17  */
  assign opb_x = n12641; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:78:10  */
  assign addsub_res = n12644; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:79:10  */
  assign cp_res = n12718; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:83:10  */
  assign cp_result = n12797; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:84:10  */
  assign cp_valid = n12798; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:85:10  */
  assign cp_shamt = n12721; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:97:10  */
  assign csr_rdata_fpu = 32'b00000000000000000000000000000000; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:97:25  */
  assign csr_rdata_cfu = 32'b00000000000000000000000000000000; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:103:20  */
  assign n12610 = rs1_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:103:49  */
  assign n12611 = n12604[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:103:38  */
  assign n12612 = ~n12611;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:103:33  */
  assign n12613 = n12610 & n12612;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:103:64  */
  assign n12614 = {n12613, rs1_i};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:104:20  */
  assign n12615 = rs2_i[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:104:49  */
  assign n12616 = n12604[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:104:38  */
  assign n12617 = ~n12616;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:104:33  */
  assign n12618 = n12615 & n12617;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:104:64  */
  assign n12619 = {n12618, rs2_i};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:106:39  */
  assign n12621 = rs1_i == rs2_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:106:27  */
  assign n12622 = n12621 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:107:49  */
  assign n12625 = $signed(cmp_rs1) < $signed(cmp_rs2);
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:107:27  */
  assign n12626 = n12625 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:113:29  */
  assign n12628 = n12604[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:113:16  */
  assign n12629 = n12628 ? pc_i : rs1_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:114:29  */
  assign n12630 = n12604[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:114:16  */
  assign n12631 = n12630 ? imm_i : rs2_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:119:16  */
  assign n12632 = opa[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:119:43  */
  assign n12633 = n12604[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:119:32  */
  assign n12634 = ~n12633;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:119:27  */
  assign n12635 = n12632 & n12634;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:119:58  */
  assign n12636 = {n12635, opa};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:120:16  */
  assign n12637 = opb[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:120:43  */
  assign n12638 = n12604[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:120:32  */
  assign n12639 = ~n12638;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:120:27  */
  assign n12640 = n12637 & n12639;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:120:58  */
  assign n12641 = {n12640, opb};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:122:51  */
  assign n12642 = opa_x - opb_x;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:122:83  */
  assign n12643 = n12604[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:122:70  */
  assign n12644 = n12643 ? n12642 : n12645;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:123:51  */
  assign n12645 = opa_x + opb_x;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:125:22  */
  assign n12646 = addsub_res[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:133:17  */
  assign n12648 = n12604[20:18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:134:7  */
  assign n12650 = n12648 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:135:48  */
  assign n12651 = addsub_res[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:135:7  */
  assign n12653 = n12648 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:136:7  */
  assign n12655 = n12648 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:137:51  */
  assign n12656 = addsub_res[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:137:7  */
  assign n12658 = n12648 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:138:7  */
  assign n12660 = n12648 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:139:42  */
  assign n12661 = opb ^ rs1_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:139:7  */
  assign n12663 = n12648 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:140:42  */
  assign n12664 = opb | rs1_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:140:7  */
  assign n12666 = n12648 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:141:42  */
  assign n12667 = opb & rs1_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:141:7  */
  assign n12669 = n12648 == 3'b111;
  assign n12670 = {n12669, n12666, n12663, n12660, n12658, n12655, n12653, n12650};
  assign n12672 = n12651[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12673 = cp_res[0]; // extract
  assign n12674 = opb[0]; // extract
  assign n12675 = n12661[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:107:7  */
  assign n12676 = n12664[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1016:3  */
  assign n12677 = n12667[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:133:5  */
  always @*
    case (n12670)
      8'b10000000: n12679 = n12677;
      8'b01000000: n12679 = n12676;
      8'b00100000: n12679 = n12675;
      8'b00010000: n12679 = n12674;
      8'b00001000: n12679 = n12656;
      8'b00000100: n12679 = n12673;
      8'b00000010: n12679 = n12672;
      8'b00000001: n12679 = 1'b0;
      default: n12679 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:107:7  */
  assign n12681 = n12651[31:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1152:14  */
  assign n12682 = cp_res[31:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12683 = opb[31:1]; // extract
  assign n12684 = n12661[31:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1253:65  */
  assign n12685 = n12664[31:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:107:7  */
  assign n12686 = n12667[31:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:133:5  */
  always @*
    case (n12670)
      8'b10000000: n12689 = n12686;
      8'b01000000: n12689 = n12685;
      8'b00100000: n12689 = n12684;
      8'b00010000: n12689 = n12683;
      8'b00001000: n12689 = 31'b0000000000000000000000000000000;
      8'b00000100: n12689 = n12682;
      8'b00000010: n12689 = n12681;
      8'b00000001: n12689 = 31'b0000000000000000000000000000000;
      default: n12689 = 31'b0000000000000000000000000000000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:24  */
  assign n12693 = cp_valid[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:39  */
  assign n12694 = cp_valid[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:28  */
  assign n12695 = n12693 | n12694;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:54  */
  assign n12696 = cp_valid[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:43  */
  assign n12697 = n12695 | n12696;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:69  */
  assign n12698 = cp_valid[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:58  */
  assign n12699 = n12697 | n12698;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:84  */
  assign n12700 = cp_valid[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:73  */
  assign n12701 = n12699 | n12700;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:99  */
  assign n12702 = cp_valid[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:88  */
  assign n12703 = n12701 | n12702;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:114  */
  assign n12704 = cp_valid[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:153:103  */
  assign n12705 = n12703 | n12704;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:22  */
  assign n12706 = cp_result[223:192]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:38  */
  assign n12707 = cp_result[191:160]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:26  */
  assign n12708 = n12706 | n12707;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:54  */
  assign n12709 = cp_result[159:128]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:42  */
  assign n12710 = n12708 | n12709;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:70  */
  assign n12711 = cp_result[127:96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:58  */
  assign n12712 = n12710 | n12711;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:86  */
  assign n12713 = cp_result[95:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:74  */
  assign n12714 = n12712 | n12713;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:102  */
  assign n12715 = cp_result[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:90  */
  assign n12716 = n12714 | n12715;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:118  */
  assign n12717 = cp_result[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:157:106  */
  assign n12718 = n12716 | n12717;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:161:32  */
  assign n12719 = csr_rdata_fpu | csr_rdata_cfu;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:164:18  */
  assign n12721 = opb[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:169:3  */
  neorv32_cpu_cp_shifter_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_cpu_cp_shifter_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .\ctrl_i_ctrl_i[if_fence] (n12722),
    .\ctrl_i_ctrl_i[rf_wb_en] (n12723),
    .\ctrl_i_ctrl_i[rf_rs1] (n12724),
    .\ctrl_i_ctrl_i[rf_rs2] (n12725),
    .\ctrl_i_ctrl_i[rf_rd] (n12726),
    .\ctrl_i_ctrl_i[rf_zero_we] (n12727),
    .\ctrl_i_ctrl_i[alu_op] (n12728),
    .\ctrl_i_ctrl_i[alu_sub] (n12729),
    .\ctrl_i_ctrl_i[alu_opa_mux] (n12730),
    .\ctrl_i_ctrl_i[alu_opb_mux] (n12731),
    .\ctrl_i_ctrl_i[alu_unsigned] (n12732),
    .\ctrl_i_ctrl_i[alu_cp_alu] (n12733),
    .\ctrl_i_ctrl_i[alu_cp_cfu] (n12734),
    .\ctrl_i_ctrl_i[alu_cp_fpu] (n12735),
    .\ctrl_i_ctrl_i[lsu_req] (n12736),
    .\ctrl_i_ctrl_i[lsu_rw] (n12737),
    .\ctrl_i_ctrl_i[lsu_mo_we] (n12738),
    .\ctrl_i_ctrl_i[lsu_fence] (n12739),
    .\ctrl_i_ctrl_i[lsu_priv] (n12740),
    .\ctrl_i_ctrl_i[ir_funct3] (n12741),
    .\ctrl_i_ctrl_i[ir_funct12] (n12742),
    .\ctrl_i_ctrl_i[ir_opcode] (n12743),
    .\ctrl_i_ctrl_i[cpu_priv] (n12744),
    .\ctrl_i_ctrl_i[cpu_sleep] (n12745),
    .\ctrl_i_ctrl_i[cpu_trap] (n12746),
    .\ctrl_i_ctrl_i[cpu_debug] (n12747),
    .rs1_i(rs1_i),
    .shamt_i(cp_shamt),
    .res_o(\neorv32_cpu_cp_shifter_inst.res_o ),
    .valid_o(\neorv32_cpu_cp_shifter_inst.valid_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:711:12  */
  assign n12722 = n12604[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12723 = n12604[1]; // extract
  assign n12724 = n12604[6:2]; // extract
  assign n12725 = n12604[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:107:7  */
  assign n12726 = n12604[16:12]; // extract
  assign n12727 = n12604[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12728 = n12604[20:18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:711:12  */
  assign n12729 = n12604[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:711:12  */
  assign n12730 = n12604[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:107:7  */
  assign n12731 = n12604[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1026:14  */
  assign n12732 = n12604[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12733 = n12604[25]; // extract
  assign n12734 = n12604[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:711:12  */
  assign n12735 = n12604[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:107:7  */
  assign n12736 = n12604[28]; // extract
  assign n12737 = n12604[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12738 = n12604[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:711:12  */
  assign n12739 = n12604[31]; // extract
  assign n12740 = n12604[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:107:7  */
  assign n12741 = n12604[35:33]; // extract
  assign n12742 = n12604[47:36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12743 = n12604[54:48]; // extract
  assign n12744 = n12604[55]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2128:5  */
  assign n12745 = n12604[56]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:107:7  */
  assign n12746 = n12604[57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:65:10  */
  assign n12747 = n12604[58]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_alu.vhd:191:5  */
  neorv32_cpu_cp_muldiv_3f29546453678b855931c174a97d6c0894b8f546 neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .\ctrl_i_ctrl_i[if_fence] (n12750),
    .\ctrl_i_ctrl_i[rf_wb_en] (n12751),
    .\ctrl_i_ctrl_i[rf_rs1] (n12752),
    .\ctrl_i_ctrl_i[rf_rs2] (n12753),
    .\ctrl_i_ctrl_i[rf_rd] (n12754),
    .\ctrl_i_ctrl_i[rf_zero_we] (n12755),
    .\ctrl_i_ctrl_i[alu_op] (n12756),
    .\ctrl_i_ctrl_i[alu_sub] (n12757),
    .\ctrl_i_ctrl_i[alu_opa_mux] (n12758),
    .\ctrl_i_ctrl_i[alu_opb_mux] (n12759),
    .\ctrl_i_ctrl_i[alu_unsigned] (n12760),
    .\ctrl_i_ctrl_i[alu_cp_alu] (n12761),
    .\ctrl_i_ctrl_i[alu_cp_cfu] (n12762),
    .\ctrl_i_ctrl_i[alu_cp_fpu] (n12763),
    .\ctrl_i_ctrl_i[lsu_req] (n12764),
    .\ctrl_i_ctrl_i[lsu_rw] (n12765),
    .\ctrl_i_ctrl_i[lsu_mo_we] (n12766),
    .\ctrl_i_ctrl_i[lsu_fence] (n12767),
    .\ctrl_i_ctrl_i[lsu_priv] (n12768),
    .\ctrl_i_ctrl_i[ir_funct3] (n12769),
    .\ctrl_i_ctrl_i[ir_funct12] (n12770),
    .\ctrl_i_ctrl_i[ir_opcode] (n12771),
    .\ctrl_i_ctrl_i[cpu_priv] (n12772),
    .\ctrl_i_ctrl_i[cpu_sleep] (n12773),
    .\ctrl_i_ctrl_i[cpu_trap] (n12774),
    .\ctrl_i_ctrl_i[cpu_debug] (n12775),
    .rs1_i(rs1_i),
    .rs2_i(rs2_i),
    .res_o(\neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst.res_o ),
    .valid_o(\neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst.valid_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:125:7  */
  assign n12750 = n12604[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:125:7  */
  assign n12751 = n12604[1]; // extract
  assign n12752 = n12604[6:2]; // extract
  assign n12753 = n12604[11:7]; // extract
  assign n12754 = n12604[16:12]; // extract
  assign n12755 = n12604[17]; // extract
  assign n12756 = n12604[20:18]; // extract
  assign n12757 = n12604[21]; // extract
  assign n12758 = n12604[22]; // extract
  assign n12759 = n12604[23]; // extract
  assign n12760 = n12604[24]; // extract
  assign n12761 = n12604[25]; // extract
  assign n12762 = n12604[26]; // extract
  assign n12763 = n12604[27]; // extract
  assign n12764 = n12604[28]; // extract
  assign n12765 = n12604[29]; // extract
  assign n12766 = n12604[30]; // extract
  assign n12767 = n12604[31]; // extract
  assign n12768 = n12604[32]; // extract
  assign n12769 = n12604[35:33]; // extract
  assign n12770 = n12604[47:36]; // extract
  assign n12771 = n12604[54:48]; // extract
  assign n12772 = n12604[55]; // extract
  assign n12773 = n12604[56]; // extract
  assign n12774 = n12604[57]; // extract
  assign n12775 = n12604[58]; // extract
  assign n12796 = {n12626, n12622};
  assign n12797 = {\neorv32_cpu_cp_shifter_inst.res_o , \neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst.res_o , 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  assign n12798 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, \neorv32_cpu_cp_muldiv_inst_true_neorv32_cpu_cp_muldiv_inst.valid_o , \neorv32_cpu_cp_shifter_inst.valid_o };
  assign n12803 = {n12689, n12679};
endmodule

module neorv32_cpu_regfile_9508e90548b0440a4a61e5743b76c1e309b23b7f
  (input  clk_i,
   input  rstn_i,
   input  \ctrl_i_ctrl_i[if_fence] ,
   input  \ctrl_i_ctrl_i[rf_wb_en] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs1] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rs2] ,
   input  [4:0] \ctrl_i_ctrl_i[rf_rd] ,
   input  \ctrl_i_ctrl_i[rf_zero_we] ,
   input  [2:0] \ctrl_i_ctrl_i[alu_op] ,
   input  \ctrl_i_ctrl_i[alu_sub] ,
   input  \ctrl_i_ctrl_i[alu_opa_mux] ,
   input  \ctrl_i_ctrl_i[alu_opb_mux] ,
   input  \ctrl_i_ctrl_i[alu_unsigned] ,
   input  \ctrl_i_ctrl_i[alu_cp_alu] ,
   input  \ctrl_i_ctrl_i[alu_cp_cfu] ,
   input  \ctrl_i_ctrl_i[alu_cp_fpu] ,
   input  \ctrl_i_ctrl_i[lsu_req] ,
   input  \ctrl_i_ctrl_i[lsu_rw] ,
   input  \ctrl_i_ctrl_i[lsu_mo_we] ,
   input  \ctrl_i_ctrl_i[lsu_fence] ,
   input  \ctrl_i_ctrl_i[lsu_priv] ,
   input  [2:0] \ctrl_i_ctrl_i[ir_funct3] ,
   input  [11:0] \ctrl_i_ctrl_i[ir_funct12] ,
   input  [6:0] \ctrl_i_ctrl_i[ir_opcode] ,
   input  \ctrl_i_ctrl_i[cpu_priv] ,
   input  \ctrl_i_ctrl_i[cpu_sleep] ,
   input  \ctrl_i_ctrl_i[cpu_trap] ,
   input  \ctrl_i_ctrl_i[cpu_debug] ,
   input  [31:0] rd_i,
   output [31:0] rs1_o,
   output [31:0] rs2_o,
   output [31:0] rs3_o);
  wire [58:0] n12013;
  wire [1023:0] reg_file;
  wire n12018;
  wire [4:0] n12021;
  wire n12023;
  wire n12024;
  wire n12025;
  wire n12033;
  wire [4:0] n12036;
  wire n12038;
  wire n12039;
  wire n12040;
  wire n12048;
  wire [4:0] n12051;
  wire n12053;
  wire n12054;
  wire n12055;
  wire n12063;
  wire [4:0] n12066;
  wire n12068;
  wire n12069;
  wire n12070;
  wire n12078;
  wire [4:0] n12081;
  wire n12083;
  wire n12084;
  wire n12085;
  wire n12093;
  wire [4:0] n12096;
  wire n12098;
  wire n12099;
  wire n12100;
  wire n12108;
  wire [4:0] n12111;
  wire n12113;
  wire n12114;
  wire n12115;
  wire n12123;
  wire [4:0] n12126;
  wire n12128;
  wire n12129;
  wire n12130;
  wire n12138;
  wire [4:0] n12141;
  wire n12143;
  wire n12144;
  wire n12145;
  wire n12153;
  wire [4:0] n12156;
  wire n12158;
  wire n12159;
  wire n12160;
  wire n12168;
  wire [4:0] n12171;
  wire n12173;
  wire n12174;
  wire n12175;
  wire n12183;
  wire [4:0] n12186;
  wire n12188;
  wire n12189;
  wire n12190;
  wire n12198;
  wire [4:0] n12201;
  wire n12203;
  wire n12204;
  wire n12205;
  wire n12213;
  wire [4:0] n12216;
  wire n12218;
  wire n12219;
  wire n12220;
  wire n12228;
  wire [4:0] n12231;
  wire n12233;
  wire n12234;
  wire n12235;
  wire n12243;
  wire [4:0] n12246;
  wire n12248;
  wire n12249;
  wire n12250;
  wire n12258;
  wire [4:0] n12261;
  wire n12263;
  wire n12264;
  wire n12265;
  wire n12273;
  wire [4:0] n12276;
  wire n12278;
  wire n12279;
  wire n12280;
  wire n12288;
  wire [4:0] n12291;
  wire n12293;
  wire n12294;
  wire n12295;
  wire n12303;
  wire [4:0] n12306;
  wire n12308;
  wire n12309;
  wire n12310;
  wire n12318;
  wire [4:0] n12321;
  wire n12323;
  wire n12324;
  wire n12325;
  wire n12333;
  wire [4:0] n12336;
  wire n12338;
  wire n12339;
  wire n12340;
  wire n12348;
  wire [4:0] n12351;
  wire n12353;
  wire n12354;
  wire n12355;
  wire n12363;
  wire [4:0] n12366;
  wire n12368;
  wire n12369;
  wire n12370;
  wire n12378;
  wire [4:0] n12381;
  wire n12383;
  wire n12384;
  wire n12385;
  wire n12393;
  wire [4:0] n12396;
  wire n12398;
  wire n12399;
  wire n12400;
  wire n12408;
  wire [4:0] n12411;
  wire n12413;
  wire n12414;
  wire n12415;
  wire n12423;
  wire [4:0] n12426;
  wire n12428;
  wire n12429;
  wire n12430;
  wire n12438;
  wire [4:0] n12441;
  wire n12443;
  wire n12444;
  wire n12445;
  wire n12453;
  wire [4:0] n12456;
  wire n12458;
  wire n12459;
  wire n12460;
  wire n12468;
  wire [4:0] n12471;
  wire n12473;
  wire n12474;
  wire n12475;
  wire n12484;
  wire [4:0] n12486;
  wire [4:0] n12490;
  localparam [31:0] n12501 = 32'b00000000000000000000000000000000;
  wire [31:0] n12502;
  wire [31:0] n12503;
  reg [31:0] n12504;
  wire [31:0] n12505;
  wire [31:0] n12506;
  reg [31:0] n12507;
  wire [31:0] n12508;
  wire [31:0] n12509;
  reg [31:0] n12510;
  wire [31:0] n12511;
  wire [31:0] n12512;
  reg [31:0] n12513;
  wire [31:0] n12514;
  wire [31:0] n12515;
  reg [31:0] n12516;
  wire [31:0] n12517;
  wire [31:0] n12518;
  reg [31:0] n12519;
  wire [31:0] n12520;
  wire [31:0] n12521;
  reg [31:0] n12522;
  wire [31:0] n12523;
  wire [31:0] n12524;
  reg [31:0] n12525;
  wire [31:0] n12526;
  wire [31:0] n12527;
  reg [31:0] n12528;
  wire [31:0] n12529;
  wire [31:0] n12530;
  reg [31:0] n12531;
  wire [31:0] n12532;
  wire [31:0] n12533;
  reg [31:0] n12534;
  wire [31:0] n12535;
  wire [31:0] n12536;
  reg [31:0] n12537;
  wire [31:0] n12538;
  wire [31:0] n12539;
  reg [31:0] n12540;
  wire [31:0] n12541;
  wire [31:0] n12542;
  reg [31:0] n12543;
  wire [31:0] n12544;
  wire [31:0] n12545;
  reg [31:0] n12546;
  wire [31:0] n12547;
  wire [31:0] n12548;
  reg [31:0] n12549;
  wire [31:0] n12550;
  wire [31:0] n12551;
  reg [31:0] n12552;
  wire [31:0] n12553;
  wire [31:0] n12554;
  reg [31:0] n12555;
  wire [31:0] n12556;
  wire [31:0] n12557;
  reg [31:0] n12558;
  wire [31:0] n12559;
  wire [31:0] n12560;
  reg [31:0] n12561;
  wire [31:0] n12562;
  wire [31:0] n12563;
  reg [31:0] n12564;
  wire [31:0] n12565;
  wire [31:0] n12566;
  reg [31:0] n12567;
  wire [31:0] n12568;
  wire [31:0] n12569;
  reg [31:0] n12570;
  wire [31:0] n12571;
  wire [31:0] n12572;
  reg [31:0] n12573;
  wire [31:0] n12574;
  wire [31:0] n12575;
  reg [31:0] n12576;
  wire [31:0] n12577;
  wire [31:0] n12578;
  reg [31:0] n12579;
  wire [31:0] n12580;
  wire [31:0] n12581;
  reg [31:0] n12582;
  wire [31:0] n12583;
  wire [31:0] n12584;
  reg [31:0] n12585;
  wire [31:0] n12586;
  wire [31:0] n12587;
  reg [31:0] n12588;
  wire [31:0] n12589;
  wire [31:0] n12590;
  reg [31:0] n12591;
  wire [31:0] n12592;
  wire [31:0] n12593;
  reg [31:0] n12594;
  wire [1023:0] n12595;
  reg [31:0] n12600;
  reg [31:0] n12601;
  wire [31:0] n12602;
  wire [31:0] n12603;
  assign rs1_o = n12600; //(module output)
  assign rs2_o = n12601; //(module output)
  assign rs3_o = n12501; //(module output)
  assign n12013 = {\ctrl_i_ctrl_i[cpu_debug] , \ctrl_i_ctrl_i[cpu_trap] , \ctrl_i_ctrl_i[cpu_sleep] , \ctrl_i_ctrl_i[cpu_priv] , \ctrl_i_ctrl_i[ir_opcode] , \ctrl_i_ctrl_i[ir_funct12] , \ctrl_i_ctrl_i[ir_funct3] , \ctrl_i_ctrl_i[lsu_priv] , \ctrl_i_ctrl_i[lsu_fence] , \ctrl_i_ctrl_i[lsu_mo_we] , \ctrl_i_ctrl_i[lsu_rw] , \ctrl_i_ctrl_i[lsu_req] , \ctrl_i_ctrl_i[alu_cp_fpu] , \ctrl_i_ctrl_i[alu_cp_cfu] , \ctrl_i_ctrl_i[alu_cp_alu] , \ctrl_i_ctrl_i[alu_unsigned] , \ctrl_i_ctrl_i[alu_opb_mux] , \ctrl_i_ctrl_i[alu_opa_mux] , \ctrl_i_ctrl_i[alu_sub] , \ctrl_i_ctrl_i[alu_op] , \ctrl_i_ctrl_i[rf_zero_we] , \ctrl_i_ctrl_i[rf_rd] , \ctrl_i_ctrl_i[rf_rs2] , \ctrl_i_ctrl_i[rf_rs1] , \ctrl_i_ctrl_i[rf_wb_en] , \ctrl_i_ctrl_i[if_fence] };
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:59:10  */
  assign reg_file = n12595; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12018 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12021 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12023 = n12021 == 5'b00001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12024 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12025 = n12024 & n12023;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12033 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12036 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12038 = n12036 == 5'b00010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12039 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12040 = n12039 & n12038;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12048 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12051 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12053 = n12051 == 5'b00011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12054 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12055 = n12054 & n12053;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12063 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12066 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12068 = n12066 == 5'b00100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12069 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12070 = n12069 & n12068;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12078 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12081 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12083 = n12081 == 5'b00101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12084 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12085 = n12084 & n12083;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12093 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12096 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12098 = n12096 == 5'b00110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12099 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12100 = n12099 & n12098;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12108 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12111 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12113 = n12111 == 5'b00111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12114 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12115 = n12114 & n12113;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12123 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12126 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12128 = n12126 == 5'b01000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12129 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12130 = n12129 & n12128;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12138 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12141 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12143 = n12141 == 5'b01001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12144 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12145 = n12144 & n12143;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12153 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12156 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12158 = n12156 == 5'b01010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12159 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12160 = n12159 & n12158;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12168 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12171 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12173 = n12171 == 5'b01011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12174 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12175 = n12174 & n12173;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12183 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12186 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12188 = n12186 == 5'b01100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12189 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12190 = n12189 & n12188;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12198 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12201 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12203 = n12201 == 5'b01101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12204 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12205 = n12204 & n12203;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12213 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12216 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12218 = n12216 == 5'b01110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12219 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12220 = n12219 & n12218;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12228 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12231 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12233 = n12231 == 5'b01111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12234 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12235 = n12234 & n12233;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12243 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12246 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12248 = n12246 == 5'b10000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12249 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12250 = n12249 & n12248;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12258 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12261 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12263 = n12261 == 5'b10001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12264 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12265 = n12264 & n12263;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12273 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12276 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12278 = n12276 == 5'b10010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12279 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12280 = n12279 & n12278;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12288 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12291 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12293 = n12291 == 5'b10011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12294 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12295 = n12294 & n12293;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12303 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12306 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12308 = n12306 == 5'b10100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12309 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12310 = n12309 & n12308;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12318 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12321 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12323 = n12321 == 5'b10101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12324 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12325 = n12324 & n12323;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12333 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12336 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12338 = n12336 == 5'b10110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12339 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12340 = n12339 & n12338;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12348 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12351 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12353 = n12351 == 5'b10111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12354 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12355 = n12354 & n12353;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12363 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12366 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12368 = n12366 == 5'b11000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12369 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12370 = n12369 & n12368;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12378 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12381 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12383 = n12381 == 5'b11001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12384 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12385 = n12384 & n12383;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12393 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12396 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12398 = n12396 == 5'b11010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12399 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12400 = n12399 & n12398;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12408 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12411 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12413 = n12411 == 5'b11011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12414 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12415 = n12414 & n12413;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12423 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12426 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12428 = n12426 == 5'b11100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12429 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12430 = n12429 & n12428;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12438 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12441 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12443 = n12441 == 5'b11101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12444 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12445 = n12444 & n12443;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12453 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12456 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12458 = n12456 == 5'b11110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12459 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12460 = n12459 & n12458;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:20  */
  assign n12468 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:36  */
  assign n12471 = n12013[16:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:62  */
  assign n12473 = n12471 == 5'b11111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:105  */
  assign n12474 = n12013[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:112:93  */
  assign n12475 = n12474 & n12473;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:125:18  */
  assign n12484 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:129:60  */
  assign n12486 = n12013[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:130:60  */
  assign n12490 = n12013[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12502 = reg_file[1023:992]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12503 = n12475 ? rd_i : n12502;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12468)
    if (n12468)
      n12504 <= 32'b00000000000000000000000000000000;
    else
      n12504 <= n12503;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12505 = reg_file[991:960]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12506 = n12460 ? rd_i : n12505;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12453)
    if (n12453)
      n12507 <= 32'b00000000000000000000000000000000;
    else
      n12507 <= n12506;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12508 = reg_file[959:928]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12509 = n12445 ? rd_i : n12508;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12438)
    if (n12438)
      n12510 <= 32'b00000000000000000000000000000000;
    else
      n12510 <= n12509;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12511 = reg_file[927:896]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12512 = n12430 ? rd_i : n12511;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12423)
    if (n12423)
      n12513 <= 32'b00000000000000000000000000000000;
    else
      n12513 <= n12512;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12514 = reg_file[895:864]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12515 = n12415 ? rd_i : n12514;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12408)
    if (n12408)
      n12516 <= 32'b00000000000000000000000000000000;
    else
      n12516 <= n12515;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12517 = reg_file[863:832]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12518 = n12400 ? rd_i : n12517;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12393)
    if (n12393)
      n12519 <= 32'b00000000000000000000000000000000;
    else
      n12519 <= n12518;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12520 = reg_file[831:800]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12521 = n12385 ? rd_i : n12520;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12378)
    if (n12378)
      n12522 <= 32'b00000000000000000000000000000000;
    else
      n12522 <= n12521;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12523 = reg_file[799:768]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12524 = n12370 ? rd_i : n12523;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12363)
    if (n12363)
      n12525 <= 32'b00000000000000000000000000000000;
    else
      n12525 <= n12524;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12526 = reg_file[767:736]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12527 = n12355 ? rd_i : n12526;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12348)
    if (n12348)
      n12528 <= 32'b00000000000000000000000000000000;
    else
      n12528 <= n12527;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12529 = reg_file[735:704]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12530 = n12340 ? rd_i : n12529;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12333)
    if (n12333)
      n12531 <= 32'b00000000000000000000000000000000;
    else
      n12531 <= n12530;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12532 = reg_file[703:672]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12533 = n12325 ? rd_i : n12532;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12318)
    if (n12318)
      n12534 <= 32'b00000000000000000000000000000000;
    else
      n12534 <= n12533;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12535 = reg_file[671:640]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12536 = n12310 ? rd_i : n12535;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12303)
    if (n12303)
      n12537 <= 32'b00000000000000000000000000000000;
    else
      n12537 <= n12536;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12538 = reg_file[639:608]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12539 = n12295 ? rd_i : n12538;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12288)
    if (n12288)
      n12540 <= 32'b00000000000000000000000000000000;
    else
      n12540 <= n12539;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12541 = reg_file[607:576]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12542 = n12280 ? rd_i : n12541;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12273)
    if (n12273)
      n12543 <= 32'b00000000000000000000000000000000;
    else
      n12543 <= n12542;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12544 = reg_file[575:544]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12545 = n12265 ? rd_i : n12544;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12258)
    if (n12258)
      n12546 <= 32'b00000000000000000000000000000000;
    else
      n12546 <= n12545;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12547 = reg_file[543:512]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12548 = n12250 ? rd_i : n12547;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12243)
    if (n12243)
      n12549 <= 32'b00000000000000000000000000000000;
    else
      n12549 <= n12548;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12550 = reg_file[511:480]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12551 = n12235 ? rd_i : n12550;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12228)
    if (n12228)
      n12552 <= 32'b00000000000000000000000000000000;
    else
      n12552 <= n12551;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12553 = reg_file[479:448]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12554 = n12220 ? rd_i : n12553;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12213)
    if (n12213)
      n12555 <= 32'b00000000000000000000000000000000;
    else
      n12555 <= n12554;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12556 = reg_file[447:416]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12557 = n12205 ? rd_i : n12556;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12198)
    if (n12198)
      n12558 <= 32'b00000000000000000000000000000000;
    else
      n12558 <= n12557;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12559 = reg_file[415:384]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12560 = n12190 ? rd_i : n12559;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12183)
    if (n12183)
      n12561 <= 32'b00000000000000000000000000000000;
    else
      n12561 <= n12560;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12562 = reg_file[383:352]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12563 = n12175 ? rd_i : n12562;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12168)
    if (n12168)
      n12564 <= 32'b00000000000000000000000000000000;
    else
      n12564 <= n12563;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12565 = reg_file[351:320]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12566 = n12160 ? rd_i : n12565;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12153)
    if (n12153)
      n12567 <= 32'b00000000000000000000000000000000;
    else
      n12567 <= n12566;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12568 = reg_file[319:288]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12569 = n12145 ? rd_i : n12568;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12138)
    if (n12138)
      n12570 <= 32'b00000000000000000000000000000000;
    else
      n12570 <= n12569;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12571 = reg_file[287:256]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12572 = n12130 ? rd_i : n12571;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12123)
    if (n12123)
      n12573 <= 32'b00000000000000000000000000000000;
    else
      n12573 <= n12572;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12574 = reg_file[255:224]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12575 = n12115 ? rd_i : n12574;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12108)
    if (n12108)
      n12576 <= 32'b00000000000000000000000000000000;
    else
      n12576 <= n12575;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12577 = reg_file[223:192]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12578 = n12100 ? rd_i : n12577;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12093)
    if (n12093)
      n12579 <= 32'b00000000000000000000000000000000;
    else
      n12579 <= n12578;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12580 = reg_file[191:160]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12581 = n12085 ? rd_i : n12580;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12078)
    if (n12078)
      n12582 <= 32'b00000000000000000000000000000000;
    else
      n12582 <= n12581;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12583 = reg_file[159:128]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12584 = n12070 ? rd_i : n12583;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12063)
    if (n12063)
      n12585 <= 32'b00000000000000000000000000000000;
    else
      n12585 <= n12584;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12586 = reg_file[127:96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12587 = n12055 ? rd_i : n12586;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12048)
    if (n12048)
      n12588 <= 32'b00000000000000000000000000000000;
    else
      n12588 <= n12587;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12589 = reg_file[95:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12590 = n12040 ? rd_i : n12589;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12033)
    if (n12033)
      n12591 <= 32'b00000000000000000000000000000000;
    else
      n12591 <= n12590;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12592 = reg_file[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  assign n12593 = n12025 ? rd_i : n12592;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:111:9  */
  always @(posedge clk_i or posedge n12018)
    if (n12018)
      n12594 <= 32'b00000000000000000000000000000000;
    else
      n12594 <= n12593;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:109:9  */
  assign n12595 = {n12504, n12507, n12510, n12513, n12516, n12519, n12522, n12525, n12528, n12531, n12534, n12537, n12540, n12543, n12546, n12549, n12552, n12555, n12558, n12561, n12564, n12567, n12570, n12573, n12576, n12579, n12582, n12585, n12588, n12591, n12594, 32'b00000000000000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:128:7  */
  always @(posedge clk_i or posedge n12484)
    if (n12484)
      n12600 <= 32'b00000000000000000000000000000000;
    else
      n12600 <= n12602;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:128:7  */
  always @(posedge clk_i or posedge n12484)
    if (n12484)
      n12601 <= 32'b00000000000000000000000000000000;
    else
      n12601 <= n12603;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:129:27  */
  assign n12602 = reg_file[n12486 * 32 +: 32]; //(Bmux)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_regfile.vhd:130:27  */
  assign n12603 = reg_file[n12490 * 32 +: 32]; //(Bmux)
endmodule

module neorv32_cpu_control_0_1_40_d6061616ddd8e9e1dfd67ab5f4d47f4cb003c4e9
  (input  clk_i,
   input  clk_aux_i,
   input  rstn_i,
   input  [31:0] \ibus_rsp_i_ibus_rsp_i[data] ,
   input  \ibus_rsp_i_ibus_rsp_i[ack] ,
   input  \ibus_rsp_i_ibus_rsp_i[err] ,
   input  pmp_fault_i,
   input  alu_cp_done_i,
   input  [1:0] alu_cmp_i,
   input  [31:0] alu_add_i,
   input  [31:0] rf_rs1_i,
   input  [31:0] xcsr_rdata_i,
   input  irq_dbg_i,
   input  [2:0] irq_machine_i,
   input  [15:0] irq_fast_i,
   input  lsu_wait_i,
   input  [31:0] lsu_mar_i,
   input  [3:0] lsu_err_i,
   output \ctrl_o_ctrl_o[if_fence] ,
   output \ctrl_o_ctrl_o[rf_wb_en] ,
   output [4:0] \ctrl_o_ctrl_o[rf_rs1] ,
   output [4:0] \ctrl_o_ctrl_o[rf_rs2] ,
   output [4:0] \ctrl_o_ctrl_o[rf_rd] ,
   output \ctrl_o_ctrl_o[rf_zero_we] ,
   output [2:0] \ctrl_o_ctrl_o[alu_op] ,
   output \ctrl_o_ctrl_o[alu_sub] ,
   output \ctrl_o_ctrl_o[alu_opa_mux] ,
   output \ctrl_o_ctrl_o[alu_opb_mux] ,
   output \ctrl_o_ctrl_o[alu_unsigned] ,
   output \ctrl_o_ctrl_o[alu_cp_alu] ,
   output \ctrl_o_ctrl_o[alu_cp_cfu] ,
   output \ctrl_o_ctrl_o[alu_cp_fpu] ,
   output \ctrl_o_ctrl_o[lsu_req] ,
   output \ctrl_o_ctrl_o[lsu_rw] ,
   output \ctrl_o_ctrl_o[lsu_mo_we] ,
   output \ctrl_o_ctrl_o[lsu_fence] ,
   output \ctrl_o_ctrl_o[lsu_priv] ,
   output [2:0] \ctrl_o_ctrl_o[ir_funct3] ,
   output [11:0] \ctrl_o_ctrl_o[ir_funct12] ,
   output [6:0] \ctrl_o_ctrl_o[ir_opcode] ,
   output \ctrl_o_ctrl_o[cpu_priv] ,
   output \ctrl_o_ctrl_o[cpu_sleep] ,
   output \ctrl_o_ctrl_o[cpu_trap] ,
   output \ctrl_o_ctrl_o[cpu_debug] ,
   output [31:0] \ibus_req_o_ibus_req_o[addr] ,
   output [31:0] \ibus_req_o_ibus_req_o[data] ,
   output [3:0] \ibus_req_o_ibus_req_o[ben] ,
   output \ibus_req_o_ibus_req_o[stb] ,
   output \ibus_req_o_ibus_req_o[rw] ,
   output \ibus_req_o_ibus_req_o[src] ,
   output \ibus_req_o_ibus_req_o[priv] ,
   output \ibus_req_o_ibus_req_o[amo] ,
   output [3:0] \ibus_req_o_ibus_req_o[amoop] ,
   output \ibus_req_o_ibus_req_o[fence] ,
   output \ibus_req_o_ibus_req_o[sleep] ,
   output \ibus_req_o_ibus_req_o[debug] ,
   output [31:0] alu_imm_o,
   output [31:0] pc_curr_o,
   output [31:0] pc_next_o,
   output [31:0] pc_ret_o,
   output [31:0] csr_rdata_o,
   output xcsr_we_o,
   output xcsr_re_o,
   output [11:0] xcsr_addr_o,
   output [31:0] xcsr_wdata_o);
  wire n7385;
  wire n7386;
  wire [4:0] n7387;
  wire [4:0] n7388;
  wire [4:0] n7389;
  wire n7390;
  wire [2:0] n7391;
  wire n7392;
  wire n7393;
  wire n7394;
  wire n7395;
  wire n7396;
  wire n7397;
  wire n7398;
  wire n7399;
  wire n7400;
  wire n7401;
  wire n7402;
  wire n7403;
  wire [2:0] n7404;
  wire [11:0] n7405;
  wire [6:0] n7406;
  wire n7407;
  wire n7408;
  wire n7409;
  wire n7410;
  wire [31:0] n7412;
  wire [31:0] n7413;
  wire [3:0] n7414;
  wire n7415;
  wire n7416;
  wire n7417;
  wire n7418;
  wire n7419;
  wire [3:0] n7420;
  wire n7421;
  wire n7422;
  wire n7423;
  wire [33:0] n7424;
  wire [37:0] fetch_engine;
  wire [75:0] ipb;
  wire [87:0] issue_engine;
  wire [132:0] exe_engine;
  wire [132:0] exe_engine_nxt;
  wire branch_taken;
  wire [6:0] opcode;
  wire [9:0] monitor_cnt;
  wire monitor_exc;
  wire sleep_mode;
  wire [106:0] trap_ctrl;
  wire [58:0] ctrl;
  wire [58:0] ctrl_nxt;
  wire [491:0] csr;
  wire [155:0] hpmevent_cfg;
  wire [309:0] cnt;
  wire [95:0] cnt_hi_rd;
  wire [95:0] cnt_lo_rd;
  wire [11:0] cnt_event;
  wire [4:0] debug_ctrl;
  wire illegal_cmd;
  wire [2:0] csr_valid;
  wire hw_trigger_match;
  wire hw_trigger_fired;
  wire n7435;
  wire [1:0] n7441;
  wire n7442;
  wire n7443;
  wire n7444;
  wire [1:0] n7445;
  wire n7447;
  wire n7449;
  wire n7450;
  wire n7451;
  wire [1:0] n7453;
  wire [1:0] n7454;
  wire [1:0] n7455;
  wire n7457;
  wire n7458;
  wire n7459;
  wire n7460;
  wire n7461;
  wire [31:0] n7462;
  wire [31:0] n7464;
  wire [29:0] n7466;
  wire n7467;
  wire n7468;
  wire n7469;
  wire n7470;
  wire [1:0] n7473;
  wire [31:0] n7474;
  wire [1:0] n7475;
  wire [1:0] n7476;
  wire [31:0] n7477;
  wire [31:0] n7478;
  wire n7480;
  wire [30:0] n7482;
  wire [31:0] n7484;
  wire n7485;
  wire [1:0] n7487;
  reg [1:0] n7488;
  reg n7489;
  wire [31:0] n7490;
  reg [31:0] n7491;
  wire n7492;
  reg n7493;
  wire [34:0] n7494;
  wire [34:0] n7499;
  wire [29:0] n7503;
  wire [31:0] n7505;
  wire [1:0] n7507;
  wire n7509;
  wire [1:0] n7510;
  wire n7512;
  wire n7513;
  wire n7514;
  wire n7516;
  wire n7517;
  wire n7518;
  wire n7519;
  wire [15:0] n7520;
  wire [16:0] n7521;
  wire n7522;
  wire [15:0] n7523;
  wire [16:0] n7524;
  wire [1:0] n7526;
  wire n7528;
  wire n7529;
  wire n7530;
  wire n7531;
  wire n7532;
  wire n7534;
  wire n7535;
  wire n7536;
  wire [1:0] n7539;
  wire n7541;
  wire n7542;
  wire n7543;
  wire n7544;
  wire n7546;
  wire n7553;
  wire n7554;
  wire \prefetch_buffer_n1_prefetch_buffer_inst.half_o ;
  wire \prefetch_buffer_n1_prefetch_buffer_inst.free_o ;
  wire [16:0] \prefetch_buffer_n1_prefetch_buffer_inst.rdata_o ;
  wire \prefetch_buffer_n1_prefetch_buffer_inst.avail_o ;
  wire n7555;
  wire [16:0] n7556;
  wire n7557;
  wire n7559;
  wire \prefetch_buffer_n2_prefetch_buffer_inst.half_o ;
  wire \prefetch_buffer_n2_prefetch_buffer_inst.free_o ;
  wire [16:0] \prefetch_buffer_n2_prefetch_buffer_inst.rdata_o ;
  wire \prefetch_buffer_n2_prefetch_buffer_inst.avail_o ;
  wire n7562;
  wire [16:0] n7563;
  wire n7564;
  wire n7566;
  wire n7570;
  wire n7573;
  wire n7574;
  wire n7575;
  wire n7576;
  wire n7577;
  wire n7578;
  wire n7579;
  wire n7580;
  wire n7581;
  wire n7582;
  wire n7583;
  wire n7584;
  localparam [1:0] n7592 = 2'b00;
  wire n7593;
  wire n7594;
  wire [1:0] n7595;
  wire n7597;
  wire n7598;
  wire n7599;
  wire n7600;
  wire [1:0] n7602;
  wire [31:0] n7603;
  wire [33:0] n7604;
  wire n7605;
  wire n7606;
  wire n7607;
  wire n7608;
  wire n7609;
  wire n7610;
  wire [1:0] n7611;
  wire n7612;
  wire [1:0] n7614;
  wire [15:0] n7615;
  wire [17:0] n7616;
  wire [15:0] n7617;
  wire [33:0] n7618;
  wire [35:0] n7619;
  wire [34:0] n7620;
  wire n7621;
  wire [34:0] n7622;
  wire [34:0] n7623;
  wire n7624;
  wire n7625;
  wire n7626;
  wire [1:0] n7627;
  wire n7629;
  wire n7630;
  wire n7631;
  wire n7632;
  wire [1:0] n7634;
  wire [31:0] n7635;
  wire [33:0] n7636;
  wire n7637;
  wire n7638;
  wire n7639;
  wire n7640;
  wire n7641;
  wire n7642;
  wire [1:0] n7643;
  wire n7644;
  wire [1:0] n7646;
  wire [15:0] n7647;
  wire [17:0] n7648;
  wire [15:0] n7649;
  wire [33:0] n7650;
  wire [35:0] n7651;
  wire n7652;
  wire [33:0] n7653;
  wire [33:0] n7654;
  wire n7655;
  wire n7656;
  wire n7657;
  wire n7658;
  wire n7659;
  wire [35:0] n7660;
  wire [35:0] n7661;
  wire n7662;
  wire n7663;
  wire [35:0] n7664;
  wire [31:0] \issue_engine_enabled_neorv32_cpu_decompressor_inst.instr_o ;
  wire [15:0] n7666;
  wire [15:0] n7668;
  wire n7669;
  wire n7670;
  wire [15:0] n7671;
  wire [15:0] n7672;
  wire n7673;
  wire n7674;
  wire n7675;
  wire n7676;
  wire n7677;
  wire n7678;
  wire n7680;
  wire [3:0] n7682;
  wire n7684;
  wire n7685;
  wire n7687;
  wire [3:0] n7690;
  localparam [31:0] n7691 = 32'b00000000000000000000000000000000;
  wire [27:0] n7692;
  wire n7694;
  wire [3:0] n7700;
  wire [3:0] n7701;
  wire [3:0] n7702;
  wire [3:0] n7703;
  wire [3:0] n7704;
  wire [15:0] n7705;
  wire [4:0] n7706;
  wire [20:0] n7707;
  wire [5:0] n7709;
  wire [26:0] n7710;
  wire [4:0] n7711;
  wire [31:0] n7712;
  wire n7714;
  wire n7716;
  wire [3:0] n7722;
  wire [3:0] n7723;
  wire [3:0] n7724;
  wire [3:0] n7725;
  wire [3:0] n7726;
  wire [15:0] n7727;
  wire [19:0] n7728;
  wire n7730;
  wire [20:0] n7731;
  wire [5:0] n7732;
  wire [26:0] n7733;
  wire [3:0] n7734;
  wire [30:0] n7735;
  wire [31:0] n7737;
  wire n7739;
  wire [19:0] n7740;
  wire [31:0] n7742;
  wire n7744;
  wire n7746;
  wire n7747;
  wire n7749;
  wire [3:0] n7755;
  wire [3:0] n7756;
  wire [3:0] n7757;
  wire [11:0] n7758;
  wire [7:0] n7760;
  wire [19:0] n7761;
  wire n7762;
  wire [20:0] n7763;
  wire [9:0] n7764;
  wire [30:0] n7765;
  wire [31:0] n7767;
  wire n7769;
  wire n7771;
  wire n7773;
  wire [3:0] n7779;
  wire [3:0] n7780;
  wire [3:0] n7781;
  wire [3:0] n7782;
  wire [3:0] n7783;
  wire [15:0] n7784;
  wire [4:0] n7785;
  wire [20:0] n7786;
  wire [9:0] n7788;
  wire [30:0] n7789;
  wire n7790;
  wire [31:0] n7791;
  wire [4:0] n7792;
  reg [31:0] n7794;
  wire [31:0] n7795;
  wire [31:0] n7796;
  wire n7802;
  wire n7803;
  wire n7804;
  wire n7805;
  wire n7806;
  wire n7807;
  wire n7808;
  wire n7809;
  wire n7810;
  wire n7811;
  wire n7812;
  wire n7814;
  wire n7817;
  wire [132:0] n7827;
  wire [30:0] n7832;
  wire [31:0] n7834;
  wire [30:0] n7835;
  wire [31:0] n7837;
  wire [30:0] n7838;
  wire [31:0] n7840;
  wire [4:0] n7841;
  wire [6:0] n7843;
  wire [2:0] n7847;
  wire [6:0] n7848;
  wire [3:0] n7849;
  wire [31:0] n7850;
  wire n7851;
  wire [31:0] n7852;
  wire [31:0] n7853;
  wire n7866;
  wire n7867;
  wire n7868;
  wire n7869;
  localparam [58:0] n7870 = 59'b00000000000000000000000000000000000000000000000000000000000;
  wire n7875;
  wire n7877;
  wire n7878;
  wire n7880;
  wire n7881;
  reg n7883;
  wire n7888;
  wire n7890;
  wire n7891;
  wire n7893;
  wire n7894;
  wire n7896;
  wire n7897;
  wire n7899;
  wire n7900;
  wire n7902;
  wire n7903;
  wire n7905;
  wire n7906;
  wire n7908;
  wire n7909;
  wire n7911;
  wire n7912;
  reg n7914;
  wire n7915;
  wire [3:0] n7918;
  wire n7921;
  wire n7922;
  wire n7923;
  wire n7926;
  wire [30:0] n7927;
  wire [31:0] n7929;
  wire n7932;
  wire n7933;
  wire n7934;
  wire n7936;
  wire n7937;
  wire [31:0] n7938;
  wire [30:0] n7939;
  wire [31:0] n7941;
  wire n7943;
  wire [68:0] n7944;
  wire [68:0] n7945;
  wire [68:0] n7946;
  wire n7947;
  wire n7948;
  wire [3:0] n7949;
  wire [3:0] n7950;
  wire [32:0] n7951;
  wire [32:0] n7952;
  wire [32:0] n7953;
  wire [31:0] n7954;
  wire [31:0] n7955;
  wire n7956;
  wire n7957;
  wire n7958;
  wire [68:0] n7959;
  wire [3:0] n7960;
  wire [3:0] n7961;
  wire [64:0] n7962;
  wire [64:0] n7963;
  wire [64:0] n7964;
  wire n7965;
  wire n7966;
  wire n7968;
  wire n7969;
  wire n7971;
  wire n7973;
  wire n7975;
  wire n7977;
  wire n7978;
  wire n7979;
  wire [24:0] n7980;
  wire [4:0] n7981;
  wire [29:0] n7982;
  wire [31:0] n7984;
  wire [29:0] n7985;
  wire [31:0] n7987;
  wire [31:0] n7988;
  wire [31:0] n7989;
  wire [31:0] n7990;
  wire n7991;
  wire [3:0] n7994;
  wire n7995;
  wire n7997;
  wire n7998;
  wire n8000;
  wire [30:0] n8001;
  wire [31:0] n8003;
  wire [30:0] n8004;
  wire [31:0] n8006;
  wire [31:0] n8007;
  wire n8011;
  wire n8017;
  wire [30:0] n8018;
  wire [31:0] n8020;
  wire n8023;
  wire n8026;
  wire n8028;
  wire n8031;
  wire n8034;
  wire n8037;
  wire [5:0] n8039;
  reg [2:0] n8040;
  wire [1:0] n8041;
  wire n8043;
  wire n8045;
  wire n8046;
  wire n8047;
  wire n8048;
  wire n8049;
  wire n8050;
  wire n8052;
  wire n8053;
  wire n8054;
  wire n8055;
  wire n8057;
  wire n8058;
  wire n8060;
  wire n8061;
  wire n8062;
  wire n8064;
  wire n8066;
  wire n8067;
  wire n8069;
  wire n8071;
  wire n8072;
  wire n8073;
  wire n8075;
  wire n8077;
  wire n8078;
  wire n8079;
  wire n8081;
  wire n8083;
  wire n8084;
  wire n8085;
  wire n8087;
  wire n8089;
  wire n8090;
  wire n8091;
  wire n8093;
  wire n8095;
  wire n8096;
  wire n8097;
  wire n8099;
  wire n8101;
  wire n8102;
  wire n8103;
  wire n8104;
  wire n8105;
  wire [3:0] n8110;
  wire n8111;
  wire n8112;
  wire n8113;
  wire n8114;
  wire n8116;
  wire n8118;
  wire n8119;
  wire n8124;
  wire n8128;
  wire n8131;
  wire n8133;
  wire n8134;
  wire n8136;
  wire n8137;
  wire n8140;
  wire n8142;
  wire n8143;
  wire n8145;
  wire n8146;
  wire n8147;
  wire n8148;
  wire n8149;
  wire n8152;
  wire n8156;
  wire n8160;
  wire n8162;
  wire n8163;
  wire n8165;
  wire n8167;
  wire n8168;
  wire [4:0] n8169;
  wire n8171;
  wire n8172;
  wire n8175;
  wire [7:0] n8177;
  reg [3:0] n8178;
  wire n8179;
  reg n8180;
  wire n8181;
  reg n8182;
  wire [2:0] n8183;
  reg [2:0] n8184;
  wire n8185;
  reg n8186;
  wire n8187;
  reg n8188;
  wire n8189;
  reg n8190;
  wire n8191;
  reg n8192;
  wire n8193;
  reg n8194;
  reg n8195;
  wire n8197;
  wire n8199;
  wire n8200;
  wire [3:0] n8203;
  wire n8204;
  wire n8205;
  wire n8207;
  wire [30:0] n8208;
  wire [31:0] n8210;
  wire n8211;
  wire n8212;
  wire n8213;
  wire n8214;
  wire n8215;
  wire n8218;
  wire [30:0] n8220;
  wire [31:0] n8222;
  wire n8225;
  wire [3:0] n8226;
  wire [31:0] n8227;
  wire n8228;
  wire n8230;
  wire n8233;
  wire n8234;
  wire n8235;
  wire n8237;
  wire n8238;
  wire n8241;
  wire n8242;
  wire n8243;
  wire n8244;
  wire n8245;
  wire n8246;
  wire n8247;
  wire n8248;
  wire n8249;
  wire n8250;
  wire n8251;
  wire n8252;
  wire n8253;
  wire n8254;
  wire [3:0] n8256;
  wire n8257;
  wire n8258;
  wire n8260;
  wire n8261;
  wire [3:0] n8263;
  wire n8265;
  wire n8268;
  wire n8269;
  wire n8270;
  wire n8271;
  wire [2:0] n8272;
  wire n8275;
  wire n8278;
  wire n8281;
  wire n8284;
  wire [3:0] n8286;
  reg [3:0] n8287;
  reg n8288;
  reg n8289;
  wire [3:0] n8290;
  wire [1:0] n8291;
  wire [1:0] n8292;
  wire [1:0] n8293;
  wire n8295;
  wire n8297;
  wire n8298;
  wire [4:0] n8299;
  wire n8301;
  wire n8302;
  wire n8304;
  wire [10:0] n8306;
  reg n8307;
  reg n8308;
  reg [3:0] n8309;
  wire [64:0] n8310;
  reg [64:0] n8311;
  reg [31:0] n8312;
  reg [31:0] n8313;
  reg n8314;
  reg n8315;
  reg n8316;
  reg n8317;
  wire [1:0] n8318;
  reg [1:0] n8319;
  reg n8320;
  wire n8321;
  reg n8322;
  wire n8323;
  reg n8324;
  wire n8325;
  reg n8326;
  wire [2:0] n8327;
  reg [2:0] n8328;
  wire n8329;
  reg n8330;
  reg n8331;
  reg n8332;
  wire n8333;
  reg n8334;
  wire n8335;
  reg n8336;
  wire n8337;
  reg n8338;
  wire n8339;
  reg n8340;
  wire n8341;
  reg n8342;
  wire [14:0] n8346;
  wire [26:0] n8351;
  wire n8352;
  reg n8353;
  reg n8354;
  wire n8356;
  wire n8357;
  wire n8358;
  wire n8359;
  wire n8360;
  wire [4:0] n8361;
  wire [4:0] n8362;
  wire [4:0] n8363;
  wire n8364;
  wire [2:0] n8365;
  wire n8366;
  wire n8367;
  wire n8368;
  wire n8369;
  wire n8370;
  wire n8371;
  wire n8372;
  wire n8373;
  wire n8374;
  wire [3:0] n8376;
  wire n8378;
  wire n8379;
  wire n8381;
  wire n8382;
  wire n8383;
  wire n8384;
  wire n8385;
  wire [2:0] n8386;
  wire [11:0] n8387;
  wire n8388;
  wire n8389;
  wire n8390;
  wire n8392;
  wire [3:0] n8394;
  wire n8396;
  wire [9:0] n8398;
  wire [9:0] n8400;
  wire n8405;
  wire [11:0] n8408;
  wire n8412;
  wire n8414;
  wire n8415;
  wire n8417;
  wire n8418;
  wire n8420;
  wire n8421;
  wire n8425;
  wire n8427;
  wire n8428;
  wire n8430;
  wire n8431;
  wire n8434;
  wire n8436;
  wire n8437;
  wire n8439;
  wire n8440;
  wire n8442;
  wire n8443;
  wire n8445;
  wire n8446;
  wire n8448;
  wire n8449;
  wire n8451;
  wire n8452;
  wire n8454;
  wire n8455;
  wire n8457;
  wire n8458;
  wire n8460;
  wire n8461;
  wire n8463;
  wire n8464;
  wire n8466;
  wire n8467;
  wire n8469;
  wire n8470;
  wire n8472;
  wire n8473;
  wire n8475;
  wire n8476;
  wire n8478;
  wire n8479;
  wire n8481;
  wire n8482;
  wire n8484;
  wire n8485;
  wire n8487;
  wire n8488;
  wire n8490;
  wire n8491;
  wire n8495;
  wire n8497;
  wire n8498;
  wire n8500;
  wire n8501;
  wire n8505;
  wire n8507;
  wire n8508;
  wire n8510;
  wire n8511;
  wire n8513;
  wire n8514;
  wire n8516;
  wire n8517;
  wire n8519;
  wire n8520;
  wire n8522;
  wire n8523;
  wire n8525;
  wire n8526;
  wire n8528;
  wire n8529;
  wire n8531;
  wire n8532;
  wire n8534;
  wire n8535;
  wire n8537;
  wire n8538;
  wire n8540;
  wire n8541;
  wire n8543;
  wire n8544;
  wire n8546;
  wire n8547;
  wire n8549;
  wire n8550;
  wire n8552;
  wire n8553;
  wire n8555;
  wire n8556;
  wire n8558;
  wire n8559;
  wire n8561;
  wire n8562;
  wire n8566;
  wire n8568;
  wire n8569;
  wire n8571;
  wire n8572;
  wire n8574;
  wire n8575;
  wire n8577;
  wire n8578;
  wire n8580;
  wire n8581;
  wire n8583;
  wire n8584;
  wire n8586;
  wire n8587;
  wire n8589;
  wire n8590;
  wire n8592;
  wire n8593;
  wire n8595;
  wire n8596;
  wire n8598;
  wire n8599;
  wire n8601;
  wire n8602;
  wire n8604;
  wire n8605;
  wire n8607;
  wire n8608;
  wire n8610;
  wire n8611;
  wire n8613;
  wire n8614;
  wire n8616;
  wire n8617;
  wire n8619;
  wire n8620;
  wire n8622;
  wire n8623;
  wire n8625;
  wire n8626;
  wire n8628;
  wire n8629;
  wire n8631;
  wire n8632;
  wire n8634;
  wire n8635;
  wire n8637;
  wire n8638;
  wire n8640;
  wire n8641;
  wire n8643;
  wire n8644;
  wire n8646;
  wire n8647;
  wire n8649;
  wire n8650;
  wire n8652;
  wire n8653;
  wire n8655;
  wire n8656;
  wire n8658;
  wire n8659;
  wire n8661;
  wire n8662;
  wire n8664;
  wire n8665;
  wire n8667;
  wire n8668;
  wire n8670;
  wire n8671;
  wire n8673;
  wire n8674;
  wire n8676;
  wire n8677;
  wire n8679;
  wire n8680;
  wire n8684;
  wire n8686;
  wire n8687;
  wire n8689;
  wire n8690;
  wire n8692;
  wire n8693;
  wire n8695;
  wire n8696;
  wire n8698;
  wire n8699;
  wire n8701;
  wire n8702;
  wire n8704;
  wire n8705;
  wire n8709;
  wire n8711;
  wire n8712;
  wire n8714;
  wire n8715;
  wire n8719;
  wire n8721;
  wire n8722;
  wire n8724;
  wire n8725;
  wire n8727;
  wire n8728;
  wire [8:0] n8730;
  reg n8731;
  wire [1:0] n8732;
  wire n8734;
  wire [2:0] n8735;
  wire n8737;
  wire [2:0] n8738;
  wire n8740;
  wire n8741;
  wire [4:0] n8742;
  wire n8744;
  wire n8745;
  wire n8746;
  wire n8749;
  wire [7:0] n8750;
  wire n8752;
  wire n8754;
  wire n8755;
  wire n8756;
  wire n8757;
  wire n8759;
  wire n8760;
  wire n8762;
  wire [3:0] n8763;
  wire n8765;
  wire n8766;
  wire [1:0] n8767;
  wire n8769;
  wire n8770;
  wire n8771;
  wire n8772;
  wire [1:0] n8773;
  wire n8775;
  wire n8776;
  wire n8777;
  wire n8778;
  wire n8779;
  wire n8780;
  wire [1:0] n8782;
  wire n8784;
  wire n8785;
  wire n8786;
  wire n8787;
  wire n8790;
  wire n8791;
  wire n8792;
  wire [6:0] n8795;
  wire n8797;
  wire n8799;
  wire n8800;
  wire n8802;
  wire n8803;
  wire [2:0] n8804;
  wire n8806;
  wire n8809;
  wire n8811;
  wire [2:0] n8812;
  wire n8814;
  wire n8816;
  wire n8817;
  wire n8819;
  wire n8820;
  wire n8822;
  wire n8823;
  wire n8825;
  wire n8826;
  wire n8828;
  wire n8829;
  reg n8832;
  wire n8834;
  wire [2:0] n8835;
  wire n8837;
  wire n8839;
  wire n8840;
  wire n8842;
  wire n8843;
  wire n8845;
  wire n8846;
  wire n8848;
  wire n8849;
  reg n8852;
  wire n8854;
  wire [2:0] n8855;
  wire n8857;
  wire n8859;
  wire n8860;
  wire n8862;
  wire n8863;
  reg n8866;
  wire n8868;
  wire n8870;
  wire n8872;
  wire n8874;
  wire n8875;
  wire n8877;
  wire n8878;
  wire n8880;
  wire n8881;
  wire n8883;
  wire n8884;
  wire [1:0] n8885;
  wire n8887;
  wire n8890;
  wire n8892;
  wire [2:0] n8893;
  wire n8895;
  wire [4:0] n8896;
  wire n8898;
  wire [4:0] n8899;
  wire n8901;
  wire n8902;
  wire [11:0] n8903;
  wire n8905;
  wire n8907;
  wire n8908;
  wire n8909;
  wire n8910;
  wire n8911;
  wire n8913;
  wire n8914;
  wire n8915;
  wire n8917;
  wire n8918;
  wire n8919;
  wire n8920;
  wire n8921;
  wire n8923;
  wire [4:0] n8924;
  reg n8928;
  wire n8930;
  wire n8932;
  wire [2:0] n8933;
  wire n8935;
  wire n8936;
  wire n8939;
  wire n8940;
  wire n8942;
  wire [8:0] n8943;
  reg n8948;
  wire [3:0] n8952;
  wire n8954;
  wire [3:0] n8955;
  wire n8957;
  wire n8958;
  wire n8959;
  wire n8960;
  wire n8961;
  wire n8964;
  wire n8967;
  wire n8968;
  wire n8969;
  wire n8970;
  wire n8971;
  wire n8972;
  wire n8973;
  wire n8974;
  wire n8975;
  wire n8976;
  wire n8977;
  wire n8978;
  wire n8979;
  wire n8980;
  wire n8981;
  wire n8982;
  wire n8983;
  wire n8984;
  wire n8985;
  wire n8986;
  wire n8987;
  wire n8988;
  wire n8989;
  wire n8990;
  wire n8991;
  wire n8992;
  wire n8993;
  wire n8994;
  wire n8995;
  wire n8996;
  wire n8997;
  wire n8998;
  wire n8999;
  wire n9000;
  wire n9001;
  wire n9002;
  wire n9003;
  wire n9004;
  wire n9005;
  wire n9006;
  wire n9007;
  wire n9008;
  wire n9009;
  wire n9010;
  wire n9011;
  wire n9012;
  wire n9013;
  wire n9014;
  wire n9015;
  wire n9016;
  wire n9017;
  wire n9018;
  wire n9019;
  wire n9020;
  wire n9021;
  wire n9022;
  wire n9023;
  wire n9024;
  wire n9025;
  wire n9026;
  wire n9027;
  wire n9028;
  wire n9029;
  wire n9030;
  wire n9031;
  wire n9032;
  wire n9033;
  wire n9034;
  wire n9035;
  wire n9036;
  wire n9037;
  wire n9038;
  wire n9039;
  wire n9040;
  wire n9041;
  wire n9042;
  wire n9043;
  wire n9044;
  wire n9045;
  wire n9046;
  wire n9047;
  wire n9048;
  wire n9049;
  wire n9050;
  wire n9051;
  wire n9052;
  wire n9053;
  wire n9054;
  wire n9055;
  wire n9056;
  wire [10:0] n9057;
  wire n9063;
  wire n9067;
  wire n9068;
  wire n9069;
  wire n9072;
  wire n9073;
  wire n9074;
  wire n9075;
  wire n9076;
  wire n9077;
  wire n9078;
  wire n9079;
  wire n9080;
  wire n9081;
  wire n9082;
  wire n9083;
  wire n9084;
  wire n9085;
  wire n9086;
  wire n9087;
  wire n9088;
  wire n9089;
  wire n9090;
  wire n9091;
  wire n9092;
  wire n9093;
  wire n9094;
  wire n9095;
  wire n9096;
  wire n9097;
  wire n9098;
  wire n9099;
  wire n9100;
  wire n9101;
  wire n9102;
  wire n9103;
  wire n9104;
  wire n9105;
  wire n9106;
  wire n9107;
  wire n9108;
  wire n9109;
  wire n9110;
  wire n9111;
  wire n9112;
  wire n9113;
  wire n9114;
  wire n9115;
  wire n9116;
  wire n9117;
  wire n9118;
  wire n9119;
  wire n9120;
  wire n9121;
  wire n9122;
  wire n9123;
  wire n9124;
  wire n9125;
  wire n9126;
  wire n9127;
  wire n9128;
  wire n9129;
  wire n9130;
  wire n9131;
  wire n9132;
  wire n9133;
  wire n9134;
  wire n9135;
  wire n9136;
  wire n9137;
  wire n9138;
  wire n9139;
  wire n9140;
  wire n9141;
  wire n9142;
  wire n9143;
  wire n9144;
  wire n9145;
  wire n9146;
  wire n9147;
  wire n9148;
  wire n9149;
  wire n9150;
  wire n9151;
  wire n9152;
  wire n9153;
  wire n9154;
  wire n9155;
  wire n9156;
  wire n9157;
  wire n9158;
  wire n9159;
  wire n9160;
  wire n9161;
  wire n9162;
  wire n9163;
  wire n9164;
  wire n9165;
  wire n9166;
  wire n9167;
  wire n9168;
  wire n9169;
  wire n9170;
  wire n9171;
  wire n9172;
  wire n9173;
  wire n9174;
  wire n9175;
  wire n9176;
  wire n9177;
  wire n9178;
  wire n9179;
  wire n9180;
  wire n9181;
  wire n9182;
  wire n9183;
  wire n9184;
  wire n9185;
  wire n9186;
  wire n9187;
  wire n9188;
  wire n9189;
  wire n9190;
  wire n9191;
  wire n9192;
  wire n9193;
  wire n9194;
  wire n9195;
  wire n9196;
  wire n9197;
  wire n9198;
  wire n9199;
  wire n9200;
  wire n9201;
  wire n9202;
  wire n9203;
  wire n9204;
  wire n9205;
  wire n9206;
  wire n9207;
  wire n9208;
  wire n9209;
  wire n9210;
  wire n9211;
  wire n9212;
  wire n9213;
  wire n9214;
  wire [41:0] n9215;
  wire [41:0] n9218;
  wire n9222;
  wire n9226;
  wire n9228;
  wire n9230;
  wire n9232;
  wire n9234;
  wire [1:0] n9240;
  wire [6:0] n9243;
  wire n9244;
  wire n9246;
  wire n9248;
  wire n9250;
  wire n9252;
  wire n9254;
  wire n9256;
  wire n9258;
  wire n9260;
  wire n9262;
  wire n9264;
  wire n9266;
  wire n9268;
  wire n9270;
  wire n9272;
  wire n9274;
  wire n9276;
  wire n9278;
  wire n9280;
  wire n9282;
  wire n9284;
  wire n9286;
  wire n9288;
  wire n9290;
  wire n9292;
  wire n9294;
  wire n9296;
  wire n9298;
  wire [6:0] n9300;
  wire [6:0] n9301;
  wire [6:0] n9302;
  wire [6:0] n9303;
  wire [6:0] n9304;
  wire [6:0] n9305;
  wire [6:0] n9306;
  wire [6:0] n9307;
  wire [6:0] n9308;
  wire [6:0] n9309;
  wire [6:0] n9310;
  wire [6:0] n9311;
  wire [6:0] n9312;
  wire [6:0] n9313;
  wire [6:0] n9314;
  wire [6:0] n9315;
  wire [6:0] n9316;
  wire [6:0] n9317;
  wire [6:0] n9318;
  wire [6:0] n9319;
  wire [6:0] n9320;
  wire [6:0] n9321;
  wire [6:0] n9322;
  wire [6:0] n9323;
  wire [6:0] n9324;
  wire [6:0] n9325;
  wire [6:0] n9326;
  wire [6:0] n9327;
  wire [6:0] n9328;
  wire [6:0] n9329;
  wire [6:0] n9330;
  wire [6:0] n9331;
  wire [31:0] n9336;
  wire n9337;
  wire [31:0] n9338;
  wire [31:0] n9339;
  wire n9341;
  wire n9345;
  wire n9346;
  wire n9347;
  wire n9355;
  wire n9357;
  wire n9359;
  wire n9360;
  wire n9361;
  wire n9362;
  wire n9363;
  wire n9365;
  wire n9366;
  wire n9367;
  wire n9369;
  wire n9370;
  wire n9371;
  wire [3:0] n9372;
  wire n9374;
  wire n9376;
  wire n9378;
  wire n9379;
  wire n9380;
  wire n9396;
  wire n9398;
  wire n9400;
  wire n9401;
  wire n9402;
  wire n9403;
  wire n9404;
  wire n9405;
  wire n9406;
  wire n9407;
  wire n9408;
  wire n9409;
  wire n9410;
  wire n9411;
  wire n9412;
  wire n9413;
  wire n9414;
  wire n9415;
  wire n9416;
  wire n9417;
  wire n9418;
  wire n9419;
  wire n9420;
  wire [3:0] n9423;
  wire n9425;
  wire n9433;
  wire n9435;
  wire n9437;
  wire n9438;
  wire n9439;
  wire n9440;
  wire n9441;
  wire n9442;
  wire n9443;
  wire n9444;
  wire n9445;
  wire n9446;
  wire n9447;
  wire n9448;
  wire n9449;
  wire n9450;
  wire n9451;
  wire n9452;
  wire n9453;
  wire n9454;
  wire n9455;
  wire n9456;
  wire n9457;
  wire n9458;
  wire n9459;
  wire n9460;
  wire n9461;
  wire n9462;
  wire n9463;
  wire n9464;
  wire n9465;
  wire n9466;
  wire n9467;
  wire n9468;
  wire n9469;
  wire n9470;
  wire n9471;
  wire n9472;
  wire n9473;
  wire n9474;
  wire n9475;
  wire n9476;
  wire n9477;
  wire n9478;
  wire n9479;
  wire n9480;
  wire n9481;
  wire n9482;
  wire n9483;
  wire n9484;
  wire n9485;
  wire [3:0] n9488;
  wire n9490;
  wire [3:0] n9491;
  wire n9493;
  wire n9494;
  wire n9495;
  wire n9496;
  wire n9497;
  wire [3:0] n9500;
  wire n9502;
  wire n9503;
  wire [3:0] n9504;
  wire n9506;
  wire n9507;
  wire n9508;
  wire n9509;
  wire n9510;
  wire n9511;
  wire n9514;
  wire [3:0] n9516;
  wire n9518;
  wire [1:0] n9519;
  wire n9521;
  wire n9522;
  wire n9523;
  wire n9524;
  wire n9525;
  wire n9528;
  wire n9540;
  wire n9542;
  wire n9544;
  wire n9545;
  wire n9546;
  wire n9547;
  wire n9548;
  wire n9549;
  wire n9550;
  wire n9551;
  wire n9552;
  wire n9553;
  wire n9554;
  wire n9555;
  wire n9556;
  wire n9557;
  wire n9558;
  wire n9559;
  wire n9560;
  wire n9561;
  wire n9562;
  wire n9563;
  wire n9564;
  wire n9565;
  wire n9566;
  wire n9567;
  wire n9568;
  wire n9569;
  wire n9570;
  wire n9571;
  wire n9572;
  wire n9573;
  wire n9574;
  wire n9575;
  wire n9576;
  wire n9577;
  wire n9578;
  wire n9579;
  wire n9580;
  wire n9581;
  wire n9582;
  wire n9583;
  wire n9584;
  wire n9585;
  wire n9586;
  wire n9587;
  wire n9589;
  wire n9593;
  wire [11:0] n9594;
  wire n9601;
  wire n9602;
  wire [31:0] n9603;
  wire [4:0] n9604;
  wire [31:0] n9606;
  wire [1:0] n9607;
  wire [31:0] n9608;
  wire [31:0] n9609;
  wire [31:0] n9610;
  wire n9612;
  wire [31:0] n9613;
  wire [31:0] n9614;
  wire [31:0] n9615;
  wire [31:0] n9616;
  wire n9618;
  wire [31:0] n9619;
  wire [1:0] n9620;
  reg [31:0] n9621;
  wire n9622;
  wire n9623;
  wire [11:0] n9624;
  wire [31:0] n9625;
  wire n9627;
  wire n9660;
  wire n9661;
  wire n9662;
  wire n9663;
  wire n9664;
  wire [11:0] n9665;
  wire n9667;
  wire n9668;
  wire n9669;
  wire n9670;
  wire n9671;
  wire n9672;
  wire n9673;
  wire n9674;
  wire [4:0] n9675;
  wire [4:0] n9676;
  wire [4:0] n9677;
  wire [11:0] n9678;
  wire n9680;
  wire n9681;
  wire n9682;
  wire n9683;
  wire [15:0] n9684;
  wire [18:0] n9685;
  wire [18:0] n9686;
  wire [18:0] n9687;
  wire [11:0] n9688;
  wire n9690;
  wire [29:0] n9691;
  wire [30:0] n9693;
  wire n9694;
  wire [31:0] n9695;
  wire [31:0] n9696;
  wire [31:0] n9697;
  wire [11:0] n9698;
  wire n9700;
  wire n9702;
  wire n9704;
  wire n9705;
  wire n9706;
  wire [1:0] n9707;
  wire [1:0] n9708;
  wire [1:0] n9709;
  wire [11:0] n9710;
  wire n9712;
  wire [31:0] n9713;
  wire [31:0] n9714;
  wire [31:0] n9715;
  wire [11:0] n9716;
  wire n9718;
  wire [30:0] n9719;
  wire [31:0] n9721;
  wire [31:0] n9722;
  wire [31:0] n9723;
  wire [11:0] n9724;
  wire n9726;
  wire n9727;
  wire [4:0] n9728;
  wire [5:0] n9729;
  wire [5:0] n9730;
  wire [5:0] n9731;
  wire [11:0] n9732;
  wire n9734;
  wire n9735;
  wire n9736;
  wire n9737;
  wire n9738;
  wire n9739;
  wire n9740;
  wire [11:0] n9741;
  wire n9743;
  wire n9745;
  wire n9746;
  wire n9747;
  wire n9748;
  wire n9749;
  wire n9750;
  wire n9751;
  wire [3:0] n9752;
  wire [3:0] n9753;
  wire [3:0] n9754;
  wire [11:0] n9755;
  wire n9757;
  wire n9759;
  wire [30:0] n9760;
  wire [31:0] n9762;
  wire [31:0] n9763;
  wire [31:0] n9764;
  wire [11:0] n9765;
  wire n9767;
  wire n9769;
  wire [31:0] n9770;
  wire [31:0] n9771;
  wire [31:0] n9772;
  wire [11:0] n9773;
  wire n9775;
  wire n9777;
  wire n9778;
  wire n9779;
  wire n9780;
  wire n9781;
  wire n9782;
  wire n9783;
  wire [1:0] n9784;
  wire [1:0] n9785;
  wire [1:0] n9786;
  wire n9787;
  wire n9788;
  wire n9789;
  wire n9790;
  wire [2:0] n9791;
  wire [2:0] n9792;
  wire [2:0] n9793;
  wire [11:0] n9794;
  wire n9796;
  wire n9798;
  wire n9799;
  wire n9800;
  wire n9801;
  wire n9802;
  wire [30:0] n9803;
  wire [31:0] n9805;
  wire n9809;
  wire n9810;
  wire n9811;
  wire n9812;
  wire n9813;
  wire n9814;
  wire n9815;
  wire n9817;
  wire n9818;
  wire [4:0] n9819;
  wire [5:0] n9820;
  wire [30:0] n9821;
  wire [31:0] n9823;
  wire n9824;
  wire n9825;
  wire n9826;
  wire n9827;
  wire [31:0] n9829;
  wire n9830;
  wire n9831;
  wire n9833;
  wire n9835;
  wire n9837;
  wire n9838;
  wire [29:0] n9839;
  wire n9840;
  wire [31:0] n9842;
  wire [31:0] n9843;
  wire n9846;
  wire n9847;
  wire [2:0] n9848;
  wire [37:0] n9849;
  wire [63:0] n9850;
  wire [2:0] n9851;
  wire [2:0] n9852;
  wire n9853;
  wire n9854;
  wire [37:0] n9855;
  wire [37:0] n9856;
  wire [63:0] n9857;
  wire [63:0] n9858;
  wire n9859;
  wire n9861;
  wire n9862;
  wire n9863;
  wire n9864;
  wire [2:0] n9865;
  wire n9866;
  wire [30:0] n9867;
  wire [31:0] n9869;
  wire [3:0] n9870;
  wire [3:0] n9871;
  wire [3:0] n9872;
  wire [31:0] n9873;
  wire [31:0] n9874;
  wire n9875;
  wire n9876;
  wire n9878;
  wire n9879;
  wire n9880;
  wire n9882;
  wire n9884;
  wire n9885;
  wire n9886;
  wire n9888;
  wire n9890;
  wire n9892;
  wire n9893;
  wire n9894;
  wire [3:0] n9896;
  wire [2:0] n9897;
  wire [2:0] n9898;
  wire [2:0] n9899;
  wire n9900;
  wire n9901;
  wire n9902;
  wire [3:0] n9903;
  wire [3:0] n9904;
  wire [3:0] n9905;
  wire n9906;
  wire n9907;
  wire [2:0] n9908;
  wire [2:0] n9909;
  wire n9910;
  wire n9911;
  wire n9912;
  wire n9913;
  wire n9915;
  wire n9917;
  wire n9919;
  wire n9921;
  wire [3:0] n9922;
  wire [23:0] n9923;
  wire [69:0] n9924;
  wire [34:0] n9925;
  wire [66:0] n9926;
  wire [3:0] n9927;
  wire [3:0] n9928;
  wire [19:0] n9929;
  wire [19:0] n9930;
  wire [19:0] n9931;
  wire n9932;
  wire n9933;
  wire [37:0] n9934;
  wire [37:0] n9935;
  wire [31:0] n9936;
  wire [31:0] n9937;
  wire [31:0] n9938;
  wire [63:0] n9939;
  wire [63:0] n9940;
  wire [34:0] n9941;
  wire [34:0] n9942;
  wire n9944;
  wire [2:0] n9945;
  wire [2:0] n9946;
  wire [2:0] n9947;
  wire n9948;
  wire n9949;
  wire n9950;
  wire [2:0] n9951;
  wire [2:0] n9952;
  wire [2:0] n9953;
  wire [31:0] n9954;
  wire [31:0] n9955;
  wire [34:0] n9956;
  wire [34:0] n9957;
  wire [34:0] n9958;
  wire n9960;
  wire [24:0] n9963;
  wire [190:0] n9964;
  wire [66:0] n9965;
  wire [24:0] n9976;
  wire [190:0] n9977;
  wire [66:0] n9978;
  wire n9986;
  wire n9987;
  wire n9988;
  wire n9990;
  wire n9994;
  wire n9995;
  wire n9996;
  wire n9997;
  localparam [31:0] n9998 = 32'b00000000000000000000000000000000;
  wire n9999;
  wire [11:0] n10000;
  wire n10002;
  wire n10004;
  wire n10005;
  wire n10007;
  wire n10008;
  wire n10010;
  wire n10012;
  wire n10013;
  wire n10015;
  wire n10016;
  wire n10018;
  wire n10019;
  wire n10021;
  wire n10023;
  wire n10024;
  wire n10025;
  wire n10026;
  wire n10027;
  wire n10028;
  wire [1:0] n10029;
  wire n10030;
  wire n10031;
  wire n10034;
  wire n10036;
  localparam [1:0] n10050 = 2'b01;
  wire n10052;
  wire n10053;
  wire n10054;
  wire n10055;
  wire [15:0] n10056;
  wire n10058;
  wire [31:0] n10059;
  wire n10061;
  wire n10062;
  wire n10063;
  wire n10065;
  wire [31:0] n10066;
  wire n10068;
  wire [30:0] n10069;
  wire [31:0] n10071;
  wire n10073;
  wire n10074;
  wire [4:0] n10075;
  wire n10077;
  wire [31:0] n10078;
  wire n10080;
  wire n10081;
  wire n10082;
  wire n10083;
  wire [15:0] n10084;
  wire n10086;
  wire [31:0] n10087;
  wire n10089;
  wire n10091;
  wire n10093;
  wire n10094;
  wire n10096;
  wire n10097;
  wire n10099;
  wire n10100;
  wire n10102;
  wire n10103;
  wire n10105;
  wire n10106;
  wire n10108;
  wire n10109;
  wire n10111;
  wire n10112;
  wire n10114;
  wire n10115;
  wire n10117;
  wire n10118;
  wire n10120;
  wire n10121;
  wire n10123;
  wire n10124;
  wire n10126;
  wire n10127;
  wire n10129;
  wire n10130;
  wire n10132;
  wire n10133;
  wire n10135;
  wire n10136;
  wire n10138;
  wire n10139;
  wire n10141;
  wire n10142;
  wire n10144;
  wire n10145;
  wire n10147;
  wire n10148;
  wire n10149;
  wire n10150;
  wire n10152;
  wire n10154;
  wire n10156;
  wire n10158;
  wire n10160;
  wire n10162;
  wire n10164;
  wire n10166;
  wire n10168;
  wire n10170;
  wire n10172;
  wire n10174;
  wire n10176;
  wire n10178;
  wire [31:0] n10179;
  wire n10181;
  wire n10183;
  wire n10184;
  wire [31:0] n10185;
  wire n10187;
  wire n10189;
  wire n10190;
  wire n10192;
  wire n10194;
  wire n10196;
  wire n10198;
  wire n10200;
  wire n10202;
  wire n10204;
  wire n10206;
  wire n10208;
  wire n10210;
  wire n10212;
  wire n10214;
  wire n10216;
  wire [31:0] n10217;
  wire n10219;
  wire n10221;
  wire n10222;
  wire [31:0] n10223;
  wire n10225;
  wire n10227;
  wire n10228;
  wire n10230;
  wire n10232;
  wire n10234;
  wire n10236;
  wire n10238;
  wire n10240;
  wire n10242;
  wire n10244;
  wire n10246;
  wire n10248;
  wire n10250;
  wire n10252;
  wire n10254;
  localparam [31:0] n10255 = 32'b00000000000000000000000000000000;
  wire n10257;
  localparam [4:0] n10258 = 5'b10011;
  wire n10260;
  localparam [31:0] n10261 = 32'b00000001000100010000000000000000;
  wire n10263;
  localparam [9:0] n10264 = 10'b0000000000;
  wire n10266;
  wire [31:0] n10267;
  wire n10269;
  wire [31:0] n10270;
  wire n10272;
  wire [31:0] n10273;
  wire n10275;
  wire [31:0] n10276;
  wire n10278;
  wire [31:0] n10279;
  wire n10281;
  localparam [31:0] n10282 = 32'b00000001000000000000000000000110;
  wire n10284;
  wire n10347;
  wire [69:0] n10348;
  wire n10349;
  wire n10350;
  wire n10351;
  wire n10352;
  wire n10353;
  wire n10354;
  wire n10355;
  wire n10356;
  wire n10357;
  wire n10358;
  wire n10359;
  wire n10360;
  wire n10361;
  wire n10362;
  wire n10363;
  wire n10364;
  wire n10365;
  wire n10366;
  wire n10367;
  wire n10368;
  wire n10369;
  wire n10370;
  reg n10371;
  wire n10372;
  wire n10373;
  wire n10374;
  wire n10375;
  wire n10376;
  wire n10377;
  wire n10378;
  wire n10379;
  wire n10380;
  wire n10381;
  wire n10382;
  wire n10383;
  wire n10384;
  wire n10385;
  wire n10386;
  wire n10387;
  wire n10388;
  wire n10389;
  wire n10390;
  wire n10391;
  wire n10392;
  wire n10393;
  reg n10394;
  wire n10395;
  wire n10396;
  wire n10397;
  wire n10398;
  wire n10399;
  wire n10400;
  wire n10401;
  wire n10402;
  wire n10403;
  wire n10404;
  wire n10405;
  wire n10406;
  wire n10407;
  wire n10408;
  wire n10409;
  wire n10410;
  wire n10411;
  wire n10412;
  wire n10413;
  wire n10414;
  wire n10415;
  wire n10416;
  reg n10417;
  wire n10418;
  wire n10419;
  wire n10420;
  wire n10421;
  wire n10422;
  wire n10423;
  wire n10424;
  wire n10425;
  wire n10426;
  wire n10427;
  wire n10428;
  wire n10429;
  wire n10430;
  wire n10431;
  wire n10432;
  wire n10433;
  wire n10434;
  wire n10435;
  wire n10436;
  wire n10437;
  wire n10438;
  wire n10439;
  reg n10440;
  wire n10441;
  wire n10442;
  wire n10443;
  wire n10444;
  wire n10445;
  wire n10446;
  wire n10447;
  wire n10448;
  wire n10449;
  wire n10450;
  wire n10451;
  wire n10452;
  wire n10453;
  wire n10454;
  wire n10455;
  wire n10456;
  wire n10457;
  wire n10458;
  wire n10459;
  wire n10460;
  wire n10461;
  wire n10462;
  reg n10463;
  wire n10464;
  wire n10465;
  wire n10466;
  wire n10467;
  wire n10468;
  wire n10469;
  wire n10470;
  wire n10471;
  wire n10472;
  wire n10473;
  wire n10474;
  wire n10475;
  wire n10476;
  wire n10477;
  wire n10478;
  wire n10479;
  wire n10480;
  wire n10481;
  wire n10482;
  wire n10483;
  reg n10484;
  wire n10485;
  wire n10486;
  wire n10487;
  wire n10488;
  wire n10489;
  wire n10490;
  wire n10491;
  wire n10492;
  wire n10493;
  wire n10494;
  wire n10495;
  wire n10496;
  wire n10497;
  wire n10498;
  wire n10499;
  wire n10500;
  wire n10501;
  wire n10502;
  wire n10503;
  wire n10504;
  reg n10505;
  wire n10506;
  wire n10507;
  wire n10508;
  wire n10509;
  wire n10510;
  wire n10511;
  wire n10512;
  wire n10513;
  wire n10514;
  wire n10515;
  wire n10516;
  wire n10517;
  wire n10518;
  wire n10519;
  wire n10520;
  wire n10521;
  wire n10522;
  wire n10523;
  wire n10524;
  wire n10525;
  reg n10526;
  wire n10527;
  wire n10528;
  wire n10529;
  wire n10530;
  wire n10531;
  wire n10532;
  wire n10533;
  wire n10534;
  wire n10535;
  wire n10536;
  wire n10537;
  wire n10538;
  wire n10539;
  wire n10540;
  wire n10541;
  wire n10542;
  wire n10543;
  wire n10544;
  wire n10545;
  wire n10546;
  reg n10547;
  wire n10548;
  wire n10549;
  wire n10550;
  wire n10551;
  wire n10552;
  wire n10553;
  wire n10554;
  wire n10555;
  wire n10556;
  wire n10557;
  wire n10558;
  wire n10559;
  wire n10560;
  wire n10561;
  wire n10562;
  wire n10563;
  wire n10564;
  wire n10565;
  wire n10566;
  wire n10567;
  reg n10568;
  wire n10569;
  wire n10570;
  wire n10571;
  wire n10572;
  wire n10573;
  wire n10574;
  wire n10575;
  wire n10576;
  wire n10577;
  wire n10578;
  wire n10579;
  wire n10580;
  wire n10581;
  wire n10582;
  wire n10583;
  wire n10584;
  wire n10585;
  wire n10586;
  wire n10587;
  reg n10588;
  wire n10589;
  wire n10590;
  wire n10591;
  wire n10592;
  wire n10593;
  wire n10594;
  wire n10595;
  wire n10596;
  wire n10597;
  wire n10598;
  wire n10599;
  wire n10600;
  wire n10601;
  wire n10602;
  wire n10603;
  wire n10604;
  wire n10605;
  wire n10606;
  wire n10607;
  wire n10608;
  reg n10609;
  wire n10610;
  wire n10611;
  wire n10612;
  wire n10613;
  wire n10614;
  wire n10615;
  wire n10616;
  wire n10617;
  wire n10618;
  wire n10619;
  wire n10620;
  wire n10621;
  wire n10622;
  wire n10623;
  wire n10624;
  wire n10625;
  wire n10626;
  wire n10627;
  wire n10628;
  wire n10629;
  reg n10630;
  wire n10631;
  wire n10632;
  wire n10633;
  wire n10634;
  wire n10635;
  wire n10636;
  wire n10637;
  wire n10638;
  wire n10639;
  wire n10640;
  wire n10641;
  wire n10642;
  wire n10643;
  wire n10644;
  wire n10645;
  wire n10646;
  wire n10647;
  wire n10648;
  wire n10649;
  reg n10650;
  wire n10651;
  wire n10652;
  wire n10653;
  wire n10654;
  wire n10655;
  wire n10656;
  wire n10657;
  wire n10658;
  wire n10659;
  wire n10660;
  wire n10661;
  wire n10662;
  wire n10663;
  wire n10664;
  wire n10665;
  wire n10666;
  wire n10667;
  wire n10668;
  wire n10669;
  reg n10670;
  wire n10671;
  wire n10672;
  wire n10673;
  wire n10674;
  wire n10675;
  wire n10676;
  wire n10677;
  wire n10678;
  wire n10679;
  wire n10680;
  wire n10681;
  wire n10682;
  wire n10683;
  wire n10684;
  wire n10685;
  wire n10686;
  wire n10687;
  wire n10688;
  wire n10689;
  reg n10690;
  wire n10691;
  wire n10692;
  wire n10693;
  wire n10694;
  wire n10695;
  wire n10696;
  wire n10697;
  wire n10698;
  wire n10699;
  wire n10700;
  wire n10701;
  wire n10702;
  wire n10703;
  wire n10704;
  wire n10705;
  wire n10706;
  wire n10707;
  wire n10708;
  wire n10709;
  wire n10710;
  wire n10711;
  reg n10712;
  wire n10713;
  wire n10714;
  wire n10715;
  wire n10716;
  wire n10717;
  wire n10718;
  wire n10719;
  wire n10720;
  wire n10721;
  wire n10722;
  wire n10723;
  wire n10724;
  wire n10725;
  wire n10726;
  wire n10727;
  wire n10728;
  wire n10729;
  wire n10730;
  wire n10731;
  wire n10732;
  wire n10733;
  reg n10734;
  wire n10735;
  wire n10736;
  wire n10737;
  wire n10738;
  wire n10739;
  wire n10740;
  wire n10741;
  wire n10742;
  wire n10743;
  wire n10744;
  wire n10745;
  wire n10746;
  wire n10747;
  wire n10748;
  wire n10749;
  wire n10750;
  wire n10751;
  wire n10752;
  wire n10753;
  wire n10754;
  wire n10755;
  reg n10756;
  wire n10757;
  wire n10758;
  wire n10759;
  wire n10760;
  wire n10761;
  wire n10762;
  wire n10763;
  wire n10764;
  wire n10765;
  wire n10766;
  wire n10767;
  wire n10768;
  wire n10769;
  wire n10770;
  wire n10771;
  wire n10772;
  wire n10773;
  wire n10774;
  wire n10775;
  wire n10776;
  wire n10777;
  reg n10778;
  wire n10779;
  wire n10780;
  wire n10781;
  wire n10782;
  wire n10783;
  wire n10784;
  wire n10785;
  wire n10786;
  wire n10787;
  wire n10788;
  wire n10789;
  wire n10790;
  wire n10791;
  wire n10792;
  wire n10793;
  wire n10794;
  wire n10795;
  wire n10796;
  wire n10797;
  wire n10798;
  wire n10799;
  reg n10800;
  wire n10801;
  wire n10802;
  wire n10803;
  wire n10804;
  wire n10805;
  wire n10806;
  wire n10807;
  wire n10808;
  wire n10809;
  wire n10810;
  wire n10811;
  wire n10812;
  wire n10813;
  wire n10814;
  wire n10815;
  wire n10816;
  wire n10817;
  wire n10818;
  wire n10819;
  wire n10820;
  wire n10821;
  reg n10822;
  wire n10823;
  wire n10824;
  wire n10825;
  wire n10826;
  wire n10827;
  wire n10828;
  wire n10829;
  wire n10830;
  wire n10831;
  wire n10832;
  wire n10833;
  wire n10834;
  wire n10835;
  wire n10836;
  wire n10837;
  wire n10838;
  wire n10839;
  wire n10840;
  wire n10841;
  wire n10842;
  wire n10843;
  reg n10844;
  wire n10845;
  wire n10846;
  wire n10847;
  wire n10848;
  wire n10849;
  wire n10850;
  wire n10851;
  wire n10852;
  wire n10853;
  wire n10854;
  wire n10855;
  wire n10856;
  wire n10857;
  wire n10858;
  wire n10859;
  wire n10860;
  wire n10861;
  wire n10862;
  wire n10863;
  wire n10864;
  wire n10865;
  reg n10866;
  wire n10867;
  wire n10868;
  wire n10869;
  wire n10870;
  wire n10871;
  wire n10872;
  wire n10873;
  wire n10874;
  wire n10875;
  wire n10876;
  wire n10877;
  wire n10878;
  wire n10879;
  wire n10880;
  wire n10881;
  wire n10882;
  wire n10883;
  wire n10884;
  wire n10885;
  wire n10886;
  wire n10887;
  reg n10888;
  wire n10889;
  wire n10890;
  wire n10891;
  wire n10892;
  wire n10893;
  wire n10894;
  wire n10895;
  wire n10896;
  wire n10897;
  wire n10898;
  wire n10899;
  wire n10900;
  wire n10901;
  wire n10902;
  wire n10903;
  wire n10904;
  wire n10905;
  wire n10906;
  wire n10907;
  wire n10908;
  wire n10909;
  reg n10910;
  wire n10911;
  wire n10912;
  wire n10913;
  wire n10914;
  wire n10915;
  wire n10916;
  wire n10917;
  wire n10918;
  wire n10919;
  wire n10920;
  wire n10921;
  wire n10922;
  wire n10923;
  wire n10924;
  wire n10925;
  wire n10926;
  wire n10927;
  wire n10928;
  wire n10929;
  wire n10930;
  wire n10931;
  reg n10932;
  wire n10933;
  wire n10934;
  wire n10935;
  wire n10936;
  wire n10937;
  wire n10938;
  wire n10939;
  wire n10940;
  wire n10941;
  wire n10942;
  wire n10943;
  wire n10944;
  wire n10945;
  wire n10946;
  wire n10947;
  wire n10948;
  wire n10949;
  wire n10950;
  wire n10951;
  wire n10952;
  wire n10953;
  reg n10954;
  wire n10955;
  wire n10956;
  wire n10957;
  wire n10958;
  wire n10959;
  wire n10960;
  wire n10961;
  wire n10962;
  wire n10963;
  wire n10964;
  wire n10965;
  wire n10966;
  wire n10967;
  wire n10968;
  wire n10969;
  wire n10970;
  wire n10971;
  wire n10972;
  wire n10973;
  wire n10974;
  wire n10975;
  reg n10976;
  wire n10977;
  wire n10978;
  wire n10979;
  wire n10980;
  wire n10981;
  wire n10982;
  wire n10983;
  wire n10984;
  wire n10985;
  wire n10986;
  wire n10987;
  wire n10988;
  wire n10989;
  wire n10990;
  wire n10991;
  wire n10992;
  wire n10993;
  wire n10994;
  wire n10995;
  wire n10996;
  wire n10997;
  reg n10998;
  wire n10999;
  wire n11000;
  wire n11001;
  wire n11002;
  wire n11003;
  wire n11004;
  wire n11005;
  wire n11006;
  wire n11007;
  wire n11008;
  wire n11009;
  wire n11010;
  wire n11011;
  wire n11012;
  wire n11013;
  wire n11014;
  wire n11015;
  wire n11016;
  wire n11017;
  wire n11018;
  wire n11019;
  wire n11020;
  reg n11021;
  wire n11022;
  wire n11023;
  wire n11024;
  wire n11025;
  wire n11026;
  wire n11027;
  wire n11028;
  wire n11029;
  wire n11030;
  wire n11031;
  wire n11032;
  wire n11033;
  wire n11034;
  wire n11035;
  wire n11036;
  wire n11037;
  wire n11038;
  wire n11039;
  wire n11040;
  wire n11041;
  wire n11042;
  wire n11043;
  reg n11044;
  wire [31:0] n11045;
  wire [31:0] n11046;
  wire [31:0] n11054;
  wire n11056;
  wire n11061;
  wire [4:0] n11062;
  wire n11064;
  wire n11065;
  wire [3:0] n11066;
  wire n11068;
  wire n11069;
  wire [31:0] n11070;
  wire [31:0] n11071;
  wire [31:0] n11072;
  wire n11073;
  wire n11074;
  wire [4:0] n11075;
  wire n11077;
  wire n11078;
  wire [3:0] n11079;
  wire n11081;
  wire n11082;
  wire [31:0] n11083;
  wire [31:0] n11084;
  wire n11085;
  wire [31:0] n11086;
  wire [31:0] n11087;
  wire [31:0] n11088;
  wire [31:0] n11099;
  wire [32:0] n11101;
  wire n11102;
  wire [32:0] n11103;
  wire [32:0] n11104;
  wire n11106;
  wire n11111;
  wire [4:0] n11112;
  wire n11114;
  wire n11115;
  wire [3:0] n11116;
  wire n11118;
  wire n11119;
  wire [31:0] n11120;
  wire [31:0] n11121;
  wire [31:0] n11122;
  wire n11123;
  wire n11124;
  wire [4:0] n11125;
  wire n11127;
  wire n11128;
  wire [3:0] n11129;
  wire n11131;
  wire n11132;
  wire [31:0] n11133;
  wire [31:0] n11134;
  wire n11135;
  wire [31:0] n11136;
  wire [31:0] n11137;
  wire [31:0] n11138;
  wire [31:0] n11149;
  wire [32:0] n11151;
  wire n11152;
  wire [32:0] n11153;
  wire [32:0] n11154;
  wire n11156;
  wire n11161;
  wire [4:0] n11162;
  wire n11164;
  wire n11165;
  wire [3:0] n11166;
  wire n11168;
  wire n11169;
  wire [31:0] n11170;
  wire [31:0] n11171;
  wire [31:0] n11172;
  wire n11173;
  wire n11174;
  wire [4:0] n11175;
  wire n11177;
  wire n11178;
  wire [3:0] n11179;
  wire n11181;
  wire n11182;
  wire [31:0] n11183;
  wire [31:0] n11184;
  wire n11185;
  wire [31:0] n11186;
  wire [31:0] n11187;
  wire [31:0] n11188;
  wire [31:0] n11199;
  wire [32:0] n11201;
  wire n11202;
  wire [32:0] n11203;
  wire [32:0] n11204;
  wire [31:0] n11206;
  localparam [95:0] n11207 = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n11209;
  localparam [95:0] n11210 = 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [31:0] n11212;
  wire [31:0] n11213;
  wire [31:0] n11214;
  wire [31:0] n11215;
  wire n11220;
  wire n11223;
  wire n11224;
  wire n11225;
  wire n11226;
  wire n11227;
  wire n11228;
  wire n11229;
  wire n11231;
  wire n11232;
  wire n11233;
  wire n11234;
  wire n11235;
  wire n11236;
  wire n11237;
  wire [11:0] n11239;
  wire [11:0] n11240;
  wire n11246;
  wire n11248;
  wire n11250;
  wire n11251;
  wire n11252;
  wire n11253;
  wire n11254;
  wire n11255;
  wire n11256;
  wire n11257;
  wire n11258;
  wire n11259;
  wire n11260;
  wire n11261;
  wire n11262;
  wire n11263;
  wire n11264;
  wire n11265;
  wire n11266;
  wire n11267;
  wire n11268;
  wire n11269;
  wire n11270;
  wire n11271;
  wire n11272;
  wire n11273;
  wire n11274;
  wire n11275;
  wire n11276;
  wire n11277;
  wire [11:0] n11279;
  wire [11:0] n11280;
  wire n11286;
  wire n11288;
  wire n11290;
  wire n11291;
  wire n11292;
  wire n11293;
  wire n11294;
  wire n11295;
  wire n11296;
  wire n11297;
  wire n11298;
  wire n11299;
  wire n11300;
  wire n11301;
  wire n11302;
  wire n11303;
  wire n11304;
  wire n11305;
  wire n11306;
  wire n11307;
  wire n11308;
  wire n11309;
  wire n11310;
  wire n11311;
  wire n11312;
  wire n11313;
  wire n11314;
  wire n11315;
  wire n11316;
  wire n11317;
  wire [11:0] n11319;
  wire [11:0] n11320;
  wire n11326;
  wire n11328;
  wire n11330;
  wire n11331;
  wire n11332;
  wire n11333;
  wire n11334;
  wire n11335;
  wire n11336;
  wire n11337;
  wire n11338;
  wire n11339;
  wire n11340;
  wire n11341;
  wire n11342;
  wire n11343;
  wire n11344;
  wire n11345;
  wire n11346;
  wire n11347;
  wire n11348;
  wire n11349;
  wire n11350;
  wire n11351;
  wire n11352;
  wire n11353;
  wire n11354;
  wire n11355;
  wire n11356;
  wire n11357;
  wire [11:0] n11359;
  wire [11:0] n11360;
  wire n11366;
  wire n11368;
  wire n11370;
  wire n11371;
  wire n11372;
  wire n11373;
  wire n11374;
  wire n11375;
  wire n11376;
  wire n11377;
  wire n11378;
  wire n11379;
  wire n11380;
  wire n11381;
  wire n11382;
  wire n11383;
  wire n11384;
  wire n11385;
  wire n11386;
  wire n11387;
  wire n11388;
  wire n11389;
  wire n11390;
  wire n11391;
  wire n11392;
  wire n11393;
  wire n11394;
  wire n11395;
  wire n11396;
  wire n11397;
  wire [11:0] n11399;
  wire [11:0] n11400;
  wire n11406;
  wire n11408;
  wire n11410;
  wire n11411;
  wire n11412;
  wire n11413;
  wire n11414;
  wire n11415;
  wire n11416;
  wire n11417;
  wire n11418;
  wire n11419;
  wire n11420;
  wire n11421;
  wire n11422;
  wire n11423;
  wire n11424;
  wire n11425;
  wire n11426;
  wire n11427;
  wire n11428;
  wire n11429;
  wire n11430;
  wire n11431;
  wire n11432;
  wire n11433;
  wire n11434;
  wire n11435;
  wire n11436;
  wire n11437;
  wire [11:0] n11439;
  wire [11:0] n11440;
  wire n11446;
  wire n11448;
  wire n11450;
  wire n11451;
  wire n11452;
  wire n11453;
  wire n11454;
  wire n11455;
  wire n11456;
  wire n11457;
  wire n11458;
  wire n11459;
  wire n11460;
  wire n11461;
  wire n11462;
  wire n11463;
  wire n11464;
  wire n11465;
  wire n11466;
  wire n11467;
  wire n11468;
  wire n11469;
  wire n11470;
  wire n11471;
  wire n11472;
  wire n11473;
  wire n11474;
  wire n11475;
  wire n11476;
  wire n11477;
  wire [11:0] n11479;
  wire [11:0] n11480;
  wire n11486;
  wire n11488;
  wire n11490;
  wire n11491;
  wire n11492;
  wire n11493;
  wire n11494;
  wire n11495;
  wire n11496;
  wire n11497;
  wire n11498;
  wire n11499;
  wire n11500;
  wire n11501;
  wire n11502;
  wire n11503;
  wire n11504;
  wire n11505;
  wire n11506;
  wire n11507;
  wire n11508;
  wire n11509;
  wire n11510;
  wire n11511;
  wire n11512;
  wire n11513;
  wire n11514;
  wire n11515;
  wire n11516;
  wire n11517;
  wire [11:0] n11519;
  wire [11:0] n11520;
  wire n11526;
  wire n11528;
  wire n11530;
  wire n11531;
  wire n11532;
  wire n11533;
  wire n11534;
  wire n11535;
  wire n11536;
  wire n11537;
  wire n11538;
  wire n11539;
  wire n11540;
  wire n11541;
  wire n11542;
  wire n11543;
  wire n11544;
  wire n11545;
  wire n11546;
  wire n11547;
  wire n11548;
  wire n11549;
  wire n11550;
  wire n11551;
  wire n11552;
  wire n11553;
  wire n11554;
  wire n11555;
  wire n11556;
  wire n11557;
  wire [11:0] n11559;
  wire [11:0] n11560;
  wire n11566;
  wire n11568;
  wire n11570;
  wire n11571;
  wire n11572;
  wire n11573;
  wire n11574;
  wire n11575;
  wire n11576;
  wire n11577;
  wire n11578;
  wire n11579;
  wire n11580;
  wire n11581;
  wire n11582;
  wire n11583;
  wire n11584;
  wire n11585;
  wire n11586;
  wire n11587;
  wire n11588;
  wire n11589;
  wire n11590;
  wire n11591;
  wire n11592;
  wire n11593;
  wire n11594;
  wire n11595;
  wire n11596;
  wire n11597;
  wire [11:0] n11599;
  wire [11:0] n11600;
  wire n11606;
  wire n11608;
  wire n11610;
  wire n11611;
  wire n11612;
  wire n11613;
  wire n11614;
  wire n11615;
  wire n11616;
  wire n11617;
  wire n11618;
  wire n11619;
  wire n11620;
  wire n11621;
  wire n11622;
  wire n11623;
  wire n11624;
  wire n11625;
  wire n11626;
  wire n11627;
  wire n11628;
  wire n11629;
  wire n11630;
  wire n11631;
  wire n11632;
  wire n11633;
  wire n11634;
  wire n11635;
  wire n11636;
  wire n11637;
  wire [11:0] n11639;
  wire [11:0] n11640;
  wire n11646;
  wire n11648;
  wire n11650;
  wire n11651;
  wire n11652;
  wire n11653;
  wire n11654;
  wire n11655;
  wire n11656;
  wire n11657;
  wire n11658;
  wire n11659;
  wire n11660;
  wire n11661;
  wire n11662;
  wire n11663;
  wire n11664;
  wire n11665;
  wire n11666;
  wire n11667;
  wire n11668;
  wire n11669;
  wire n11670;
  wire n11671;
  wire n11672;
  wire n11673;
  wire n11674;
  wire n11675;
  wire n11676;
  wire n11677;
  wire [11:0] n11679;
  wire [11:0] n11680;
  wire n11686;
  wire n11688;
  wire n11690;
  wire n11691;
  wire n11692;
  wire n11693;
  wire n11694;
  wire n11695;
  wire n11696;
  wire n11697;
  wire n11698;
  wire n11699;
  wire n11700;
  wire n11701;
  wire n11702;
  wire n11703;
  wire n11704;
  wire n11705;
  wire n11706;
  wire n11707;
  wire n11708;
  wire n11709;
  wire n11710;
  wire n11711;
  wire n11712;
  wire n11713;
  wire n11714;
  wire n11715;
  wire n11716;
  wire n11717;
  wire [11:0] n11719;
  wire [11:0] n11720;
  wire n11726;
  wire n11728;
  wire n11730;
  wire n11731;
  wire n11732;
  wire n11733;
  wire n11734;
  wire n11735;
  wire n11736;
  wire n11737;
  wire n11738;
  wire n11739;
  wire n11740;
  wire n11741;
  wire n11742;
  wire n11743;
  wire n11744;
  wire n11745;
  wire n11746;
  wire n11747;
  wire n11748;
  wire n11749;
  wire n11750;
  wire n11751;
  wire n11752;
  wire n11753;
  wire n11754;
  wire n11755;
  wire n11756;
  wire n11757;
  wire [15:0] n11758;
  wire n11764;
  wire n11765;
  wire [3:0] n11769;
  wire n11771;
  wire n11772;
  wire [3:0] n11775;
  wire n11777;
  wire n11778;
  wire n11779;
  wire n11780;
  wire [3:0] n11783;
  wire n11785;
  wire [1:0] n11786;
  wire n11788;
  wire n11789;
  wire n11790;
  wire [3:0] n11793;
  wire n11795;
  wire n11796;
  wire [3:0] n11799;
  wire n11801;
  wire n11802;
  wire [3:0] n11805;
  wire n11807;
  wire n11808;
  wire n11811;
  wire n11812;
  wire n11813;
  wire n11814;
  wire n11815;
  wire n11816;
  wire n11817;
  wire n11820;
  wire n11821;
  wire n11822;
  wire n11823;
  wire n11824;
  wire n11825;
  wire n11828;
  wire n11829;
  wire [3:0] n11830;
  wire n11832;
  wire n11833;
  wire n11834;
  wire n11837;
  wire n11838;
  wire n11841;
  wire n11844;
  wire n11845;
  wire n11846;
  wire n11847;
  wire n11848;
  wire n11850;
  wire n11851;
  wire n11852;
  wire n11854;
  wire n11855;
  wire n11856;
  wire n11861;
  wire n11862;
  wire n11863;
  wire n11864;
  wire n11865;
  wire n11866;
  wire n11867;
  wire n11868;
  wire n11869;
  wire n11870;
  wire n11871;
  wire n11872;
  wire n11873;
  wire n11874;
  wire n11875;
  wire n11876;
  wire n11877;
  wire n11878;
  wire n11879;
  wire n11880;
  wire n11881;
  wire n11882;
  wire n11883;
  wire n11884;
  wire n11885;
  wire n11886;
  wire n11887;
  wire n11890;
  wire n11893;
  wire n11895;
  wire [2:0] n11900;
  wire n11904;
  wire n11905;
  wire n11906;
  wire [1:0] n11907;
  wire n11909;
  wire n11910;
  wire n11911;
  wire [30:0] n11912;
  wire [30:0] n11913;
  wire n11914;
  wire n11915;
  wire n11916;
  wire n11919;
  wire n11921;
  wire n11922;
  wire n11923;
  wire n11924;
  wire [11:0] n11925;
  wire n11927;
  wire n11928;
  wire n11929;
  wire n11930;
  wire n11931;
  wire n11933;
  wire n11934;
  wire n11940;
  wire n11948;
  wire [3:0] n11950;
  wire n11958;
  reg n11961;
  reg [34:0] n11962;
  wire [37:0] n11963;
  wire [75:0] n11964;
  reg n11965;
  wire [87:0] n11966;
  reg [132:0] n11967;
  wire [132:0] n11968;
  reg [9:0] n11969;
  reg n11970;
  reg n11971;
  reg n11972;
  reg [6:0] n11973;
  reg [41:0] n11974;
  reg [10:0] n11975;
  wire [106:0] n11976;
  reg [58:0] n11977;
  wire [58:0] n11978;
  reg [31:0] n11979;
  reg n11980;
  wire [31:0] n11981;
  wire [31:0] n11982;
  reg [31:0] n11983;
  reg [66:0] n11984;
  reg [190:0] n11985;
  reg [24:0] n11986;
  reg n11987;
  wire [11:0] n11988;
  wire [11:0] n11989;
  reg [11:0] n11990;
  wire [491:0] n11991;
  reg [15:0] n11992;
  reg n11993;
  reg [31:0] n11994;
  reg [31:0] n11995;
  reg n11996;
  reg [31:0] n11997;
  reg [31:0] n11998;
  reg n11999;
  reg [31:0] n12000;
  reg [31:0] n12001;
  wire [309:0] n12002;
  wire [95:0] n12003;
  wire [95:0] n12004;
  wire [11:0] n12005;
  reg n12006;
  wire [4:0] n12007;
  wire [2:0] n12008;
  reg n12009;
  wire [58:0] n12010;
  wire [79:0] n12011;
  reg [31:0] n12012;
  assign \ctrl_o_ctrl_o[if_fence]  = n7385; //(module output)
  assign \ctrl_o_ctrl_o[rf_wb_en]  = n7386; //(module output)
  assign \ctrl_o_ctrl_o[rf_rs1]  = n7387; //(module output)
  assign \ctrl_o_ctrl_o[rf_rs2]  = n7388; //(module output)
  assign \ctrl_o_ctrl_o[rf_rd]  = n7389; //(module output)
  assign \ctrl_o_ctrl_o[rf_zero_we]  = n7390; //(module output)
  assign \ctrl_o_ctrl_o[alu_op]  = n7391; //(module output)
  assign \ctrl_o_ctrl_o[alu_sub]  = n7392; //(module output)
  assign \ctrl_o_ctrl_o[alu_opa_mux]  = n7393; //(module output)
  assign \ctrl_o_ctrl_o[alu_opb_mux]  = n7394; //(module output)
  assign \ctrl_o_ctrl_o[alu_unsigned]  = n7395; //(module output)
  assign \ctrl_o_ctrl_o[alu_cp_alu]  = n7396; //(module output)
  assign \ctrl_o_ctrl_o[alu_cp_cfu]  = n7397; //(module output)
  assign \ctrl_o_ctrl_o[alu_cp_fpu]  = n7398; //(module output)
  assign \ctrl_o_ctrl_o[lsu_req]  = n7399; //(module output)
  assign \ctrl_o_ctrl_o[lsu_rw]  = n7400; //(module output)
  assign \ctrl_o_ctrl_o[lsu_mo_we]  = n7401; //(module output)
  assign \ctrl_o_ctrl_o[lsu_fence]  = n7402; //(module output)
  assign \ctrl_o_ctrl_o[lsu_priv]  = n7403; //(module output)
  assign \ctrl_o_ctrl_o[ir_funct3]  = n7404; //(module output)
  assign \ctrl_o_ctrl_o[ir_funct12]  = n7405; //(module output)
  assign \ctrl_o_ctrl_o[ir_opcode]  = n7406; //(module output)
  assign \ctrl_o_ctrl_o[cpu_priv]  = n7407; //(module output)
  assign \ctrl_o_ctrl_o[cpu_sleep]  = n7408; //(module output)
  assign \ctrl_o_ctrl_o[cpu_trap]  = n7409; //(module output)
  assign \ctrl_o_ctrl_o[cpu_debug]  = n7410; //(module output)
  assign \ibus_req_o_ibus_req_o[addr]  = n7412; //(module output)
  assign \ibus_req_o_ibus_req_o[data]  = n7413; //(module output)
  assign \ibus_req_o_ibus_req_o[ben]  = n7414; //(module output)
  assign \ibus_req_o_ibus_req_o[stb]  = n7415; //(module output)
  assign \ibus_req_o_ibus_req_o[rw]  = n7416; //(module output)
  assign \ibus_req_o_ibus_req_o[src]  = n7417; //(module output)
  assign \ibus_req_o_ibus_req_o[priv]  = n7418; //(module output)
  assign \ibus_req_o_ibus_req_o[amo]  = n7419; //(module output)
  assign \ibus_req_o_ibus_req_o[amoop]  = n7420; //(module output)
  assign \ibus_req_o_ibus_req_o[fence]  = n7421; //(module output)
  assign \ibus_req_o_ibus_req_o[sleep]  = n7422; //(module output)
  assign \ibus_req_o_ibus_req_o[debug]  = n7423; //(module output)
  assign alu_imm_o = n12012; //(module output)
  assign pc_curr_o = n7834; //(module output)
  assign pc_next_o = n7837; //(module output)
  assign pc_ret_o = n7840; //(module output)
  assign csr_rdata_o = n11054; //(module output)
  assign xcsr_we_o = n9622; //(module output)
  assign xcsr_re_o = n9623; //(module output)
  assign xcsr_addr_o = n9624; //(module output)
  assign xcsr_wdata_o = n9625; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:692:41  */
  assign n7385 = n12010[0]; // extract
  assign n7386 = n12010[1]; // extract
  assign n7387 = n12010[6:2]; // extract
  assign n7388 = n12010[11:7]; // extract
  assign n7389 = n12010[16:12]; // extract
  assign n7390 = n12010[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1038:14  */
  assign n7391 = n12010[20:18]; // extract
  assign n7392 = n12010[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n7393 = n12010[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n7394 = n12010[23]; // extract
  assign n7395 = n12010[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n7396 = n12010[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:710:68  */
  assign n7397 = n12010[26]; // extract
  assign n7398 = n12010[27]; // extract
  assign n7399 = n12010[28]; // extract
  assign n7400 = n12010[29]; // extract
  assign n7401 = n12010[30]; // extract
  assign n7402 = n12010[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:694:43  */
  assign n7403 = n12010[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:692:42  */
  assign n7404 = n12010[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:650:3  */
  assign n7405 = n12010[47:36]; // extract
  assign n7406 = n12010[54:48]; // extract
  assign n7407 = n12010[55]; // extract
  assign n7408 = n12010[56]; // extract
  assign n7409 = n12010[57]; // extract
  assign n7410 = n12010[58]; // extract
  assign n7412 = n12011[31:0]; // extract
  assign n7413 = n12011[63:32]; // extract
  assign n7414 = n12011[67:64]; // extract
  assign n7415 = n12011[68]; // extract
  assign n7416 = n12011[69]; // extract
  assign n7417 = n12011[70]; // extract
  assign n7418 = n12011[71]; // extract
  assign n7419 = n12011[72]; // extract
  assign n7420 = n12011[76:73]; // extract
  assign n7421 = n12011[77]; // extract
  assign n7422 = n12011[78]; // extract
  assign n7423 = n12011[79]; // extract
  assign n7424 = {\ibus_rsp_i_ibus_rsp_i[err] , \ibus_rsp_i_ibus_rsp_i[ack] , \ibus_rsp_i_ibus_rsp_i[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:131:10  */
  assign fetch_engine = n11963; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:140:10  */
  assign ipb = n11964; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:153:10  */
  assign issue_engine = n11966; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:166:10  */
  assign exe_engine = n11967; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:166:22  */
  assign exe_engine_nxt = n11968; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:169:10  */
  assign branch_taken = n7814; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:172:10  */
  assign opcode = n7843; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:175:10  */
  assign monitor_cnt = n11969; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:176:10  */
  assign monitor_exc = n8405; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:179:10  */
  assign sleep_mode = n11970; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:204:10  */
  assign trap_ctrl = n11976; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:207:10  */
  assign ctrl = n11977; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:207:16  */
  assign ctrl_nxt = n11978; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:257:10  */
  assign csr = n11991; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:262:10  */
  assign hpmevent_cfg = 156'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:277:10  */
  assign cnt = n12002; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:278:10  */
  assign cnt_hi_rd = n12003; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:278:21  */
  assign cnt_lo_rd = n12004; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:281:10  */
  assign cnt_event = n12005; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:287:10  */
  assign debug_ctrl = n12007; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:290:10  */
  assign illegal_cmd = n8948; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:293:10  */
  assign csr_valid = n12008; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:296:10  */
  assign hw_trigger_match = n11916; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:296:28  */
  assign hw_trigger_fired = n12009; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:308:16  */
  assign n7435 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:314:25  */
  assign n7441 = fetch_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:318:48  */
  assign n7442 = fetch_engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:318:72  */
  assign n7443 = fetch_engine[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:318:56  */
  assign n7444 = n7442 | n7443;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:319:19  */
  assign n7445 = ipb[73:72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:319:24  */
  assign n7447 = n7445 == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:321:31  */
  assign n7449 = fetch_engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:321:63  */
  assign n7450 = fetch_engine[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:321:46  */
  assign n7451 = n7449 | n7450;
  assign n7453 = fetch_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:321:11  */
  assign n7454 = n7451 ? 2'b00 : n7453;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:319:11  */
  assign n7455 = n7447 ? 2'b10 : n7454;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:316:9  */
  assign n7457 = n7441 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:327:48  */
  assign n7458 = fetch_engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:327:72  */
  assign n7459 = fetch_engine[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:327:56  */
  assign n7460 = n7458 | n7459;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:328:28  */
  assign n7461 = fetch_engine[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:329:75  */
  assign n7462 = fetch_engine[34:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:329:79  */
  assign n7464 = n7462 + 32'b00000000000000000000000000000100;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:711:12  */
  assign n7466 = n7464[31:2]; // extract
  assign n7467 = n7464[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:331:30  */
  assign n7468 = fetch_engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:331:62  */
  assign n7469 = fetch_engine[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:331:45  */
  assign n7470 = n7468 | n7469;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:331:13  */
  assign n7473 = n7470 ? 2'b00 : 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:395:3  */
  assign n7474 = {n7466, 1'b0, n7467};
  assign n7475 = fetch_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:328:11  */
  assign n7476 = n7461 ? n7473 : n7475;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:344:3  */
  assign n7477 = fetch_engine[34:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:328:11  */
  assign n7478 = n7461 ? n7474 : n7477;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:325:9  */
  assign n7480 = n7441 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:341:49  */
  assign n7482 = exe_engine[100:70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:341:67  */
  assign n7484 = {n7482, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:342:39  */
  assign n7485 = csr[137]; // extract
  assign n7487 = {n7480, n7457};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:314:7  */
  always @*
    case (n7487)
      2'b10: n7488 = n7476;
      2'b01: n7488 = n7455;
      default: n7488 = 2'b01;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:314:7  */
  always @*
    case (n7487)
      2'b10: n7489 = n7460;
      2'b01: n7489 = n7444;
      default: n7489 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1026:14  */
  assign n7490 = fetch_engine[34:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:314:7  */
  always @*
    case (n7487)
      2'b10: n7491 = n7478;
      2'b01: n7491 = n7490;
      default: n7491 = n7484;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:711:12  */
  assign n7492 = fetch_engine[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:314:7  */
  always @*
    case (n7487)
      2'b10: n7493 = n7492;
      2'b01: n7493 = n7492;
      default: n7493 = n7485;
    endcase
  assign n7494 = {n7491, n7489, n7488};
  assign n7499 = {32'b00000000000000000000000000000000, 1'b1, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:350:37  */
  assign n7503 = fetch_engine[34:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:350:55  */
  assign n7505 = {n7503, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:353:44  */
  assign n7507 = fetch_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:353:50  */
  assign n7509 = n7507 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:353:73  */
  assign n7510 = ipb[73:72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:353:78  */
  assign n7512 = n7510 == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:353:64  */
  assign n7513 = n7512 & n7509;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:353:25  */
  assign n7514 = n7513 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:356:35  */
  assign n7516 = n7424[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:356:53  */
  assign n7517 = n7424[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:356:39  */
  assign n7518 = n7516 | n7517;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:359:30  */
  assign n7519 = n7424[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:359:51  */
  assign n7520 = n7424[15:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:359:34  */
  assign n7521 = {n7519, n7520};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:360:30  */
  assign n7522 = n7424[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:360:51  */
  assign n7523 = n7424[31:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:360:34  */
  assign n7524 = {n7522, n7523};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:363:39  */
  assign n7526 = fetch_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:363:45  */
  assign n7528 = n7526 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:363:77  */
  assign n7529 = fetch_engine[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:363:59  */
  assign n7530 = n7529 & n7528;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:364:42  */
  assign n7531 = fetch_engine[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:364:46  */
  assign n7532 = ~n7531;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:364:53  */
  assign n7534 = n7532 | 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:363:89  */
  assign n7535 = n7534 & n7530;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:363:20  */
  assign n7536 = n7535 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:365:39  */
  assign n7539 = fetch_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:365:45  */
  assign n7541 = n7539 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:365:77  */
  assign n7542 = fetch_engine[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:365:59  */
  assign n7543 = n7542 & n7541;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:365:20  */
  assign n7544 = n7543 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:368:36  */
  assign n7546 = fetch_engine[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:375:28  */
  assign n7553 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:377:34  */
  assign n7554 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:384:5  */
  neorv32_fifo_2_17_29e2dcfbb16f63bb0254df7585a15bb6fb5e927d prefetch_buffer_n1_prefetch_buffer_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n7555),
    .wdata_i(n7556),
    .we_i(n7557),
    .re_i(n7559),
    .half_o(),
    .free_o(\prefetch_buffer_n1_prefetch_buffer_inst.free_o ),
    .rdata_o(\prefetch_buffer_n1_prefetch_buffer_inst.rdata_o ),
    .avail_o(\prefetch_buffer_n1_prefetch_buffer_inst.avail_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:396:31  */
  assign n7555 = fetch_engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:399:27  */
  assign n7556 = ipb[33:17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:400:24  */
  assign n7557 = ipb[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:403:24  */
  assign n7559 = ipb[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:384:5  */
  neorv32_fifo_2_17_29e2dcfbb16f63bb0254df7585a15bb6fb5e927d prefetch_buffer_n2_prefetch_buffer_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n7562),
    .wdata_i(n7563),
    .we_i(n7564),
    .re_i(n7566),
    .half_o(),
    .free_o(\prefetch_buffer_n2_prefetch_buffer_inst.free_o ),
    .rdata_o(\prefetch_buffer_n2_prefetch_buffer_inst.rdata_o ),
    .avail_o(\prefetch_buffer_n2_prefetch_buffer_inst.avail_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:396:31  */
  assign n7562 = fetch_engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:399:27  */
  assign n7563 = ipb[16:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:400:24  */
  assign n7564 = ipb[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:403:24  */
  assign n7566 = ipb[71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:421:18  */
  assign n7570 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:424:26  */
  assign n7573 = fetch_engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:425:47  */
  assign n7574 = exe_engine[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:426:29  */
  assign n7575 = issue_engine[87]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:427:47  */
  assign n7576 = issue_engine[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:427:75  */
  assign n7577 = issue_engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:427:58  */
  assign n7578 = ~n7577;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:427:53  */
  assign n7579 = n7576 & n7578;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:427:103  */
  assign n7580 = issue_engine[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:427:87  */
  assign n7581 = n7579 | n7580;
  assign n7582 = issue_engine[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:426:9  */
  assign n7583 = n7575 ? n7581 : n7582;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:424:9  */
  assign n7584 = n7573 ? n7574 : n7583;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:439:24  */
  assign n7593 = issue_engine[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:439:30  */
  assign n7594 = ~n7593;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:440:25  */
  assign n7595 = ipb[52:51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:440:38  */
  assign n7597 = n7595 != 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:441:46  */
  assign n7598 = ipb[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:442:46  */
  assign n7599 = ipb[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:443:55  */
  assign n7600 = ipb[67]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:443:41  */
  assign n7602 = {1'b1, n7600};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:443:75  */
  assign n7603 = issue_engine[50:19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:443:60  */
  assign n7604 = {n7602, n7603};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:445:54  */
  assign n7605 = ipb[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:445:71  */
  assign n7606 = ipb[75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:445:58  */
  assign n7607 = n7605 & n7606;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:445:54  */
  assign n7608 = ipb[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:445:71  */
  assign n7609 = ipb[75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:445:58  */
  assign n7610 = n7608 & n7609;
  assign n7611 = {n7607, n7610};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:446:51  */
  assign n7612 = ipb[67]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:446:37  */
  assign n7614 = {1'b0, n7612};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:446:70  */
  assign n7615 = ipb[49:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:446:56  */
  assign n7616 = {n7614, n7615};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:446:98  */
  assign n7617 = ipb[66:51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:446:84  */
  assign n7618 = {n7616, n7617};
  assign n7619 = {n7611, n7618};
  assign n7620 = {n7599, n7604};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:439:7  */
  assign n7621 = n7662 ? n7598 : 1'b0;
  assign n7622 = n7619[34:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:440:9  */
  assign n7623 = n7597 ? n7620 : n7622;
  assign n7624 = n7619[35]; // extract
  assign n7625 = n7592[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:440:9  */
  assign n7626 = n7597 ? n7625 : n7624;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:450:25  */
  assign n7627 = ipb[35:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:450:38  */
  assign n7629 = n7627 != 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:451:46  */
  assign n7630 = ipb[75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:452:46  */
  assign n7631 = ipb[75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:453:55  */
  assign n7632 = ipb[50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:453:41  */
  assign n7634 = {1'b1, n7632};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:453:75  */
  assign n7635 = issue_engine[50:19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:453:60  */
  assign n7636 = {n7634, n7635};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:455:54  */
  assign n7637 = ipb[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:455:71  */
  assign n7638 = ipb[75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:455:58  */
  assign n7639 = n7637 & n7638;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:455:54  */
  assign n7640 = ipb[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:455:71  */
  assign n7641 = ipb[75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:455:58  */
  assign n7642 = n7640 & n7641;
  assign n7643 = {n7639, n7642};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:456:51  */
  assign n7644 = ipb[67]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:456:37  */
  assign n7646 = {1'b0, n7644};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:456:70  */
  assign n7647 = ipb[66:51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:456:56  */
  assign n7648 = {n7646, n7647};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:456:98  */
  assign n7649 = ipb[49:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:456:84  */
  assign n7650 = {n7648, n7649};
  assign n7651 = {n7643, n7650};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:450:9  */
  assign n7652 = n7629 ? n7630 : 1'b0;
  assign n7653 = n7651[33:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:450:9  */
  assign n7654 = n7629 ? n7636 : n7653;
  assign n7655 = n7651[34]; // extract
  assign n7656 = n7592[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:450:9  */
  assign n7657 = n7629 ? n7656 : n7655;
  assign n7658 = n7651[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:450:9  */
  assign n7659 = n7629 ? n7631 : n7658;
  assign n7660 = {n7659, n7657, n7654};
  assign n7661 = {n7626, n7623};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:439:7  */
  assign n7662 = n7597 & n7594;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:439:7  */
  assign n7663 = n7594 ? 1'b0 : n7652;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:439:7  */
  assign n7664 = n7594 ? n7661 : n7660;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:464:5  */
  neorv32_cpu_decompressor issue_engine_enabled_neorv32_cpu_decompressor_inst (
    .instr_i(n7666),
    .instr_o(\issue_engine_enabled_neorv32_cpu_decompressor_inst.instr_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:466:31  */
  assign n7666 = issue_engine[18:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:471:40  */
  assign n7668 = ipb[66:51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:471:73  */
  assign n7669 = issue_engine[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:471:79  */
  assign n7670 = ~n7669;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:471:54  */
  assign n7671 = n7670 ? n7668 : n7672;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:471:103  */
  assign n7672 = ipb[49:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:489:34  */
  assign n7673 = issue_engine[85]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:489:55  */
  assign n7674 = issue_engine[87]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:489:38  */
  assign n7675 = n7673 & n7674;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:490:34  */
  assign n7676 = issue_engine[86]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:490:55  */
  assign n7677 = issue_engine[87]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:490:38  */
  assign n7678 = n7676 & n7677;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:501:16  */
  assign n7680 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:504:22  */
  assign n7682 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:504:28  */
  assign n7684 = n7682 == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:506:46  */
  assign n7685 = issue_engine[84]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:506:24  */
  assign n7687 = n7685 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:506:9  */
  assign n7690 = n7687 ? 4'b0010 : 4'b0100;
  assign n7692 = n7691[31:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:514:51  */
  assign n7694 = exe_engine[35]; // extract
  assign n7700 = {n7694, n7694, n7694, n7694};
  assign n7701 = {n7694, n7694, n7694, n7694};
  assign n7702 = {n7694, n7694, n7694, n7694};
  assign n7703 = {n7694, n7694, n7694, n7694};
  assign n7704 = {n7694, n7694, n7694, n7694};
  assign n7705 = {n7700, n7701, n7702, n7703};
  assign n7706 = {n7704, n7694};
  assign n7707 = {n7705, n7706};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:514:76  */
  assign n7709 = exe_engine[34:29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:514:61  */
  assign n7710 = {n7707, n7709};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:514:106  */
  assign n7711 = exe_engine[15:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:514:91  */
  assign n7712 = {n7710, n7711};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:513:11  */
  assign n7714 = opcode == 7'b0100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:516:51  */
  assign n7716 = exe_engine[35]; // extract
  assign n7722 = {n7716, n7716, n7716, n7716};
  assign n7723 = {n7716, n7716, n7716, n7716};
  assign n7724 = {n7716, n7716, n7716, n7716};
  assign n7725 = {n7716, n7716, n7716, n7716};
  assign n7726 = {n7716, n7716, n7716, n7716};
  assign n7727 = {n7722, n7723, n7724, n7725};
  assign n7728 = {n7727, n7726};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:516:76  */
  assign n7730 = exe_engine[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:516:61  */
  assign n7731 = {n7728, n7730};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:516:95  */
  assign n7732 = exe_engine[34:29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:516:80  */
  assign n7733 = {n7731, n7732};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:516:125  */
  assign n7734 = exe_engine[15:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:516:110  */
  assign n7735 = {n7733, n7734};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:516:139  */
  assign n7737 = {n7735, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:515:11  */
  assign n7739 = opcode == 7'b1100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:518:39  */
  assign n7740 = exe_engine[35:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:518:54  */
  assign n7742 = {n7740, 12'b000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:517:11  */
  assign n7744 = opcode == 7'b0110111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:517:29  */
  assign n7746 = opcode == 7'b0010111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:517:29  */
  assign n7747 = n7744 | n7746;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:520:51  */
  assign n7749 = exe_engine[35]; // extract
  assign n7755 = {n7749, n7749, n7749, n7749};
  assign n7756 = {n7749, n7749, n7749, n7749};
  assign n7757 = {n7749, n7749, n7749, n7749};
  assign n7758 = {n7755, n7756, n7757};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:520:76  */
  assign n7760 = exe_engine[23:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:520:61  */
  assign n7761 = {n7758, n7760};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:520:106  */
  assign n7762 = exe_engine[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:520:91  */
  assign n7763 = {n7761, n7762};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:520:126  */
  assign n7764 = exe_engine[34:25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:520:111  */
  assign n7765 = {n7763, n7764};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:520:141  */
  assign n7767 = {n7765, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:519:11  */
  assign n7769 = opcode == 7'b1101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:521:11  */
  assign n7771 = opcode == 7'b0101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:524:51  */
  assign n7773 = exe_engine[35]; // extract
  assign n7779 = {n7773, n7773, n7773, n7773};
  assign n7780 = {n7773, n7773, n7773, n7773};
  assign n7781 = {n7773, n7773, n7773, n7773};
  assign n7782 = {n7773, n7773, n7773, n7773};
  assign n7783 = {n7773, n7773, n7773, n7773};
  assign n7784 = {n7779, n7780, n7781, n7782};
  assign n7785 = {n7783, n7773};
  assign n7786 = {n7784, n7785};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:524:76  */
  assign n7788 = exe_engine[34:25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:524:61  */
  assign n7789 = {n7786, n7788};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:524:106  */
  assign n7790 = exe_engine[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:524:91  */
  assign n7791 = {n7789, n7790};
  assign n7792 = {n7771, n7769, n7747, n7739, n7714};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:512:9  */
  always @*
    case (n7792)
      5'b10000: n7794 = 32'b00000000000000000000000000000000;
      5'b01000: n7794 = n7767;
      5'b00100: n7794 = n7742;
      5'b00010: n7794 = n7737;
      5'b00001: n7794 = n7712;
      default: n7794 = n7791;
    endcase
  assign n7795 = {n7692, n7690};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:504:7  */
  assign n7796 = n7684 ? n7795 : n7794;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:535:22  */
  assign n7802 = exe_engine[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:535:45  */
  assign n7803 = ~n7802;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:536:24  */
  assign n7804 = exe_engine[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:536:45  */
  assign n7805 = ~n7804;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:537:34  */
  assign n7806 = alu_cmp_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:537:65  */
  assign n7807 = exe_engine[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:537:48  */
  assign n7808 = n7806 ^ n7807;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:539:34  */
  assign n7809 = alu_cmp_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:539:64  */
  assign n7810 = exe_engine[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:539:47  */
  assign n7811 = n7809 ^ n7810;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:536:7  */
  assign n7812 = n7805 ? n7808 : n7811;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:535:5  */
  assign n7814 = n7803 ? n7812 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:551:16  */
  assign n7817 = ~rstn_i;
  assign n7827 = {32'b00000000000000000000000000000000, 32'b11111111111000000000000000000000, 32'b11111111111000000000000000000000, 1'b0, 32'b00000000000000000000000000000000, 4'b0011};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:566:29  */
  assign n7832 = exe_engine[68:38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:566:47  */
  assign n7834 = {n7832, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:567:30  */
  assign n7835 = exe_engine[100:70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:567:48  */
  assign n7837 = {n7835, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:568:29  */
  assign n7838 = exe_engine[132:102]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:568:47  */
  assign n7840 = {n7838, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:571:26  */
  assign n7841 = exe_engine[10:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:571:75  */
  assign n7843 = {n7841, 2'b11};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:582:30  */
  assign n7847 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:583:30  */
  assign n7848 = exe_engine[35:29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:586:40  */
  assign n7849 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:587:40  */
  assign n7850 = exe_engine[35:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:588:40  */
  assign n7851 = exe_engine[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:589:40  */
  assign n7852 = exe_engine[68:37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:590:40  */
  assign n7853 = exe_engine[100:69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:606:15  */
  assign n7866 = opcode[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:607:40  */
  assign n7867 = exe_engine[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:609:40  */
  assign n7868 = exe_engine[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:606:5  */
  assign n7869 = n7866 ? n7867 : n7868;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:614:7  */
  assign n7875 = opcode == 7'b0010111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:614:27  */
  assign n7877 = opcode == 7'b1101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:614:27  */
  assign n7878 = n7875 | n7877;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:614:42  */
  assign n7880 = opcode == 7'b1100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:614:42  */
  assign n7881 = n7878 | n7880;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:613:5  */
  always @*
    case (n7881)
      1'b1: n7883 = 1'b1;
      default: n7883 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:7  */
  assign n7888 = opcode == 7'b0010011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:26  */
  assign n7890 = opcode == 7'b0110111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:26  */
  assign n7891 = n7888 | n7890;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:41  */
  assign n7893 = opcode == 7'b0010111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:41  */
  assign n7894 = n7891 | n7893;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:58  */
  assign n7896 = opcode == 7'b0000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:58  */
  assign n7897 = n7894 | n7896;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:74  */
  assign n7899 = opcode == 7'b0100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:74  */
  assign n7900 = n7897 | n7899;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:91  */
  assign n7902 = opcode == 7'b0101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:91  */
  assign n7903 = n7900 | n7902;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:106  */
  assign n7905 = opcode == 7'b1100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:106  */
  assign n7906 = n7903 | n7905;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:124  */
  assign n7908 = opcode == 7'b1101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:124  */
  assign n7909 = n7906 | n7908;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:139  */
  assign n7911 = opcode == 7'b1100111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:622:139  */
  assign n7912 = n7909 | n7911;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:621:5  */
  always @*
    case (n7912)
      1'b1: n7914 = 1'b1;
      default: n7914 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:632:39  */
  assign n7915 = exe_engine[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:21  */
  assign n7918 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:643:23  */
  assign n7921 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:643:56  */
  assign n7922 = trap_ctrl[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:643:42  */
  assign n7923 = n7921 | n7922;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:645:32  */
  assign n7926 = hw_trigger_match & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:646:49  */
  assign n7927 = exe_engine[100:70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:646:67  */
  assign n7929 = {n7927, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:649:34  */
  assign n7932 = issue_engine[85]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:649:67  */
  assign n7933 = issue_engine[86]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:649:45  */
  assign n7934 = n7932 | n7933;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:651:52  */
  assign n7936 = issue_engine[83]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:652:52  */
  assign n7937 = issue_engine[84]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:653:52  */
  assign n7938 = issue_engine[82:51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:654:49  */
  assign n7939 = exe_engine[100:70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:654:67  */
  assign n7941 = {n7939, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:649:9  */
  assign n7943 = n7934 ? 1'b1 : 1'b0;
  assign n7944 = {n7941, n7937, n7938, 4'b0101};
  assign n7945 = {n7852, n7851, n7850, n7849};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:649:9  */
  assign n7946 = n7934 ? n7944 : n7945;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:649:9  */
  assign n7947 = n7934 ? n7936 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:645:9  */
  assign n7948 = n7926 ? 1'b0 : n7943;
  assign n7949 = n7946[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:645:9  */
  assign n7950 = n7926 ? 4'b0000 : n7949;
  assign n7951 = n7946[36:4]; // extract
  assign n7952 = {n7851, n7850};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:645:9  */
  assign n7953 = n7926 ? n7952 : n7951;
  assign n7954 = n7946[68:37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:645:9  */
  assign n7955 = n7926 ? n7929 : n7954;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:645:9  */
  assign n7956 = n7926 ? 1'b0 : n7947;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:645:9  */
  assign n7957 = n7926 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:643:9  */
  assign n7958 = n7923 ? 1'b0 : n7948;
  assign n7959 = {n7955, n7953, n7950};
  assign n7960 = n7959[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:643:9  */
  assign n7961 = n7923 ? 4'b0001 : n7960;
  assign n7962 = n7959[68:4]; // extract
  assign n7963 = {n7852, n7851, n7850};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:643:9  */
  assign n7964 = n7923 ? n7963 : n7962;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:643:9  */
  assign n7965 = n7923 ? 1'b0 : n7956;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:643:9  */
  assign n7966 = n7923 ? 1'b0 : n7957;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:638:7  */
  assign n7968 = n7918 == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:660:28  */
  assign n7969 = trap_ctrl[62]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:660:39  */
  assign n7971 = 1'b1 & n7969;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:662:27  */
  assign n7973 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:662:38  */
  assign n7975 = 1'b1 & n7973;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:665:24  */
  assign n7977 = csr[176]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:665:55  */
  assign n7978 = trap_ctrl[63]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:665:35  */
  assign n7979 = n7978 & n7977;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:666:44  */
  assign n7980 = csr[207:183]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:666:79  */
  assign n7981 = trap_ctrl[61:57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:666:62  */
  assign n7982 = {n7980, n7981};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:666:92  */
  assign n7984 = {n7982, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:668:44  */
  assign n7985 = csr[207:178]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:668:62  */
  assign n7987 = {n7985, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:665:11  */
  assign n7988 = n7979 ? n7984 : n7987;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:662:9  */
  assign n7989 = n7975 ? 32'b11111111111111111111111000000000 : n7988;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:660:9  */
  assign n7990 = n7971 ? 32'b11111111111111111111111000010000 : n7989;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:672:23  */
  assign n7991 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:672:9  */
  assign n7994 = n7991 ? 4'b0011 : n7849;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:672:9  */
  assign n7995 = n7991 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:658:7  */
  assign n7997 = n7918 == 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:679:24  */
  assign n7998 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:679:35  */
  assign n8000 = 1'b1 & n7998;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:680:40  */
  assign n8001 = csr[392:362]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:680:58  */
  assign n8003 = {n8001, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:682:41  */
  assign n8004 = csr[169:139]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:682:59  */
  assign n8006 = {n8004, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:679:9  */
  assign n8007 = n8000 ? n8003 : n8006;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:677:7  */
  assign n8011 = n7918 == 4'b0010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:687:7  */
  assign n8017 = n7918 == 4'b0011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:695:40  */
  assign n8018 = alu_add_i[31:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:695:58  */
  assign n8020 = {n8018, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:706:15  */
  assign n8023 = n7847 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:707:15  */
  assign n8026 = n7847 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:708:15  */
  assign n8028 = n7847 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:709:15  */
  assign n8031 = n7847 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:710:15  */
  assign n8034 = n7847 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:711:15  */
  assign n8037 = n7847 == 3'b111;
  assign n8039 = {n8037, n8034, n8031, n8028, n8026, n8023};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:705:13  */
  always @*
    case (n8039)
      6'b100000: n8040 = 3'b111;
      6'b010000: n8040 = 3'b110;
      6'b001000: n8040 = 3'b101;
      6'b000100: n8040 = 3'b011;
      6'b000010: n8040 = 3'b011;
      6'b000001: n8040 = 3'b001;
      default: n8040 = 3'b000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:716:25  */
  assign n8041 = exe_engine[18:17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:716:38  */
  assign n8043 = n8041 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:717:27  */
  assign n8045 = n7847 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:717:55  */
  assign n8046 = opcode[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:717:44  */
  assign n8047 = n8046 & n8045;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:717:84  */
  assign n8048 = exe_engine[34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:717:66  */
  assign n8049 = n8048 & n8047;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:716:66  */
  assign n8050 = n8043 | n8049;
  assign n8052 = n7870[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:716:13  */
  assign n8053 = n8050 ? 1'b1 : n8052;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:24  */
  assign n8054 = opcode[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:28  */
  assign n8055 = ~n8054;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:49  */
  assign n8057 = n7847 != 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:35  */
  assign n8058 = n8057 & n8055;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:80  */
  assign n8060 = n7847 != 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:66  */
  assign n8061 = n8060 & n8058;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:24  */
  assign n8062 = opcode[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:51  */
  assign n8064 = n7847 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:82  */
  assign n8066 = n7848 == 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:68  */
  assign n8067 = n8066 & n8064;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:110  */
  assign n8069 = n7847 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:141  */
  assign n8071 = n7848 == 7'b0100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:127  */
  assign n8072 = n8071 & n8069;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:96  */
  assign n8073 = n8067 | n8072;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:724:51  */
  assign n8075 = n7847 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:724:82  */
  assign n8077 = n7848 == 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:724:68  */
  assign n8078 = n8077 & n8075;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:155  */
  assign n8079 = n8073 | n8078;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:724:110  */
  assign n8081 = n7847 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:724:141  */
  assign n8083 = n7848 == 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:724:127  */
  assign n8084 = n8083 & n8081;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:724:96  */
  assign n8085 = n8079 | n8084;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:725:51  */
  assign n8087 = n7847 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:725:82  */
  assign n8089 = n7848 == 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:725:68  */
  assign n8090 = n8089 & n8087;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:724:155  */
  assign n8091 = n8085 | n8090;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:725:110  */
  assign n8093 = n7847 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:725:141  */
  assign n8095 = n7848 == 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:725:127  */
  assign n8096 = n8095 & n8093;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:725:96  */
  assign n8097 = n8091 | n8096;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:726:51  */
  assign n8099 = n7847 == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:726:82  */
  assign n8101 = n7848 == 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:726:68  */
  assign n8102 = n8101 & n8099;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:725:155  */
  assign n8103 = n8097 | n8102;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:723:35  */
  assign n8104 = n8103 & n8062;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:97  */
  assign n8105 = n8061 | n8104;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:13  */
  assign n8110 = n8105 ? 4'b0000 : 4'b0110;
  assign n8111 = n7870[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:13  */
  assign n8112 = n8105 ? 1'b1 : n8111;
  assign n8113 = n7870[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:722:13  */
  assign n8114 = n8105 ? n8113 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:702:11  */
  assign n8116 = opcode == 7'b0110011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:702:29  */
  assign n8118 = opcode == 7'b0010011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:702:29  */
  assign n8119 = n8116 | n8118;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:735:11  */
  assign n8124 = opcode == 7'b0110111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:741:11  */
  assign n8128 = opcode == 7'b0010111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:747:11  */
  assign n8131 = opcode == 7'b0000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:747:30  */
  assign n8133 = opcode == 7'b0100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:747:30  */
  assign n8134 = n8131 | n8133;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:747:47  */
  assign n8136 = opcode == 7'b0101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:747:47  */
  assign n8137 = n8134 | n8136;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:751:11  */
  assign n8140 = opcode == 7'b1100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:751:32  */
  assign n8142 = opcode == 7'b1101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:751:32  */
  assign n8143 = n8140 | n8142;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:751:47  */
  assign n8145 = opcode == 7'b1100111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:751:47  */
  assign n8146 = n8143 | n8145;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:756:54  */
  assign n8147 = exe_engine[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:757:54  */
  assign n8148 = exe_engine[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:757:37  */
  assign n8149 = ~n8148;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:755:11  */
  assign n8152 = opcode == 7'b0001111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:761:11  */
  assign n8156 = opcode == 7'b1010011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:766:11  */
  assign n8160 = opcode == 7'b0001011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:766:31  */
  assign n8162 = opcode == 7'b0101011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:766:31  */
  assign n8163 = n8160 | n8162;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:772:27  */
  assign n8165 = n7847 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:772:58  */
  assign n8167 = n7847 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:772:45  */
  assign n8168 = n8165 | n8167;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:772:96  */
  assign n8169 = exe_engine[15:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:772:135  */
  assign n8171 = n8169 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:772:78  */
  assign n8172 = n8171 & n8168;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:772:13  */
  assign n8175 = n8172 ? 1'b0 : 1'b1;
  assign n8177 = {n8163, n8156, n8152, n8146, n8137, n8128, n8124, n8119};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8178 = 4'b0110;
      8'b01000000: n8178 = 4'b0110;
      8'b00100000: n8178 = 4'b0011;
      8'b00010000: n8178 = 4'b0111;
      8'b00001000: n8178 = 4'b1010;
      8'b00000100: n8178 = 4'b0000;
      8'b00000010: n8178 = 4'b0000;
      8'b00000001: n8178 = n8110;
      default: n8178 = 4'b1001;
    endcase
  assign n8179 = n7870[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8180 = n8179;
      8'b01000000: n8180 = n8179;
      8'b00100000: n8180 = n8147;
      8'b00010000: n8180 = n8179;
      8'b00001000: n8180 = n8179;
      8'b00000100: n8180 = n8179;
      8'b00000010: n8180 = n8179;
      8'b00000001: n8180 = n8179;
      default: n8180 = n8179;
    endcase
  assign n8181 = n7870[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8182 = n8181;
      8'b01000000: n8182 = n8181;
      8'b00100000: n8182 = n8181;
      8'b00010000: n8182 = n8181;
      8'b00001000: n8182 = n8181;
      8'b00000100: n8182 = 1'b1;
      8'b00000010: n8182 = 1'b1;
      8'b00000001: n8182 = n8112;
      default: n8182 = n8181;
    endcase
  assign n8183 = n7870[20:18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8184 = n8183;
      8'b01000000: n8184 = n8183;
      8'b00100000: n8184 = n8183;
      8'b00010000: n8184 = n8183;
      8'b00001000: n8184 = n8183;
      8'b00000100: n8184 = 3'b001;
      8'b00000010: n8184 = 3'b100;
      8'b00000001: n8184 = n8040;
      default: n8184 = n8183;
    endcase
  assign n8185 = n7870[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8186 = n8185;
      8'b01000000: n8186 = n8185;
      8'b00100000: n8186 = n8185;
      8'b00010000: n8186 = n8185;
      8'b00001000: n8186 = n8185;
      8'b00000100: n8186 = n8185;
      8'b00000010: n8186 = n8185;
      8'b00000001: n8186 = n8053;
      default: n8186 = n8185;
    endcase
  assign n8187 = n7870[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8188 = n8187;
      8'b01000000: n8188 = n8187;
      8'b00100000: n8188 = n8187;
      8'b00010000: n8188 = n8187;
      8'b00001000: n8188 = n8187;
      8'b00000100: n8188 = n8187;
      8'b00000010: n8188 = n8187;
      8'b00000001: n8188 = n8114;
      default: n8188 = n8187;
    endcase
  assign n8189 = n7870[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8190 = 1'b1;
      8'b01000000: n8190 = n8189;
      8'b00100000: n8190 = n8189;
      8'b00010000: n8190 = n8189;
      8'b00001000: n8190 = n8189;
      8'b00000100: n8190 = n8189;
      8'b00000010: n8190 = n8189;
      8'b00000001: n8190 = n8189;
      default: n8190 = n8189;
    endcase
  assign n8191 = n7870[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8192 = n8191;
      8'b01000000: n8192 = 1'b1;
      8'b00100000: n8192 = n8191;
      8'b00010000: n8192 = n8191;
      8'b00001000: n8192 = n8191;
      8'b00000100: n8192 = n8191;
      8'b00000010: n8192 = n8191;
      8'b00000001: n8192 = n8191;
      default: n8192 = n8191;
    endcase
  assign n8193 = n7870[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8194 = n8193;
      8'b01000000: n8194 = n8193;
      8'b00100000: n8194 = n8149;
      8'b00010000: n8194 = n8193;
      8'b00001000: n8194 = n8193;
      8'b00000100: n8194 = n8193;
      8'b00000010: n8194 = n8193;
      8'b00000001: n8194 = n8193;
      default: n8194 = n8193;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:699:9  */
  always @*
    case (n8177)
      8'b10000000: n8195 = 1'b0;
      8'b01000000: n8195 = 1'b0;
      8'b00100000: n8195 = 1'b0;
      8'b00010000: n8195 = 1'b0;
      8'b00001000: n8195 = 1'b0;
      8'b00000100: n8195 = 1'b0;
      8'b00000010: n8195 = 1'b0;
      8'b00000001: n8195 = 1'b0;
      default: n8195 = n8175;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:693:7  */
  assign n8197 = n7918 == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:784:55  */
  assign n8199 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:784:34  */
  assign n8200 = alu_cp_done_i | n8199;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:784:9  */
  assign n8203 = n8200 ? 4'b0000 : n7849;
  assign n8204 = n7870[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:784:9  */
  assign n8205 = n8200 ? 1'b1 : n8204;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:781:7  */
  assign n8207 = n7918 == 4'b0110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:791:44  */
  assign n8208 = exe_engine[100:70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:791:62  */
  assign n8210 = {n8208, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:792:36  */
  assign n8211 = opcode[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:793:30  */
  assign n8212 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:793:46  */
  assign n8213 = ~n8212;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:793:53  */
  assign n8214 = branch_taken & n8213;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:794:44  */
  assign n8215 = alu_add_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:794:48  */
  assign n8218 = n8215 & 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:796:44  */
  assign n8220 = alu_add_i[31:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:796:62  */
  assign n8222 = {n8220, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:793:9  */
  assign n8225 = n8214 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:793:9  */
  assign n8226 = n8214 ? 4'b1000 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:793:9  */
  assign n8227 = n8214 ? n8222 : n7853;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:793:9  */
  assign n8228 = n8214 ? n8218 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:789:7  */
  assign n8230 = n7918 == 4'b0111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:802:7  */
  assign n8233 = n7918 == 4'b1000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:808:30  */
  assign n8234 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:808:46  */
  assign n8235 = ~n8234;
  assign n8237 = n7870[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:808:9  */
  assign n8238 = n8235 ? 1'b1 : n8237;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:806:7  */
  assign n8241 = n7918 == 4'b1010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:815:24  */
  assign n8242 = ~lsu_wait_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:816:30  */
  assign n8243 = trap_ctrl[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:815:31  */
  assign n8244 = n8242 | n8243;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:816:74  */
  assign n8245 = trap_ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:816:53  */
  assign n8246 = n8244 | n8245;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:817:30  */
  assign n8247 = trap_ctrl[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:816:97  */
  assign n8248 = n8246 | n8247;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:817:74  */
  assign n8249 = trap_ctrl[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:817:53  */
  assign n8250 = n8248 | n8249;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:818:30  */
  assign n8251 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:817:97  */
  assign n8252 = n8250 | n8251;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:819:44  */
  assign n8253 = ctrl[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:819:35  */
  assign n8254 = ~n8253;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:815:9  */
  assign n8256 = n8252 ? 4'b0000 : n7849;
  assign n8257 = n7870[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:815:9  */
  assign n8258 = n8252 ? n8254 : n8257;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:813:7  */
  assign n8260 = n7918 == 4'b1011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:825:23  */
  assign n8261 = trap_ctrl[100]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:825:9  */
  assign n8263 = n8261 ? 4'b0000 : n7849;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:823:7  */
  assign n8265 = n7918 == 4'b0100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:832:22  */
  assign n8268 = n7847 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:832:60  */
  assign n8269 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:832:76  */
  assign n8270 = ~n8269;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:832:38  */
  assign n8271 = n8270 & n8268;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:833:29  */
  assign n8272 = exe_engine[26:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:834:13  */
  assign n8275 = n8272 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:835:13  */
  assign n8278 = n8272 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:836:13  */
  assign n8281 = n8272 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:837:13  */
  assign n8284 = n8272 == 3'b101;
  assign n8286 = {n8284, n8281, n8278, n8275};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:833:11  */
  always @*
    case (n8286)
      4'b1000: n8287 = 4'b0100;
      4'b0100: n8287 = 4'b0010;
      4'b0010: n8287 = 4'b0000;
      4'b0001: n8287 = 4'b0000;
      default: n8287 = 4'b0000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:833:11  */
  always @*
    case (n8286)
      4'b1000: n8288 = 1'b0;
      4'b0100: n8288 = 1'b0;
      4'b0010: n8288 = 1'b0;
      4'b0001: n8288 = 1'b1;
      default: n8288 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:833:11  */
  always @*
    case (n8286)
      4'b1000: n8289 = 1'b0;
      4'b0100: n8289 = 1'b0;
      4'b0010: n8289 = 1'b1;
      4'b0001: n8289 = 1'b0;
      default: n8289 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:832:9  */
  assign n8290 = n8271 ? n8287 : 4'b0000;
  assign n8291 = {n8289, n8288};
  assign n8292 = {1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:832:9  */
  assign n8293 = n8271 ? n8291 : n8292;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:842:22  */
  assign n8295 = n7847 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:842:53  */
  assign n8297 = n7847 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:842:40  */
  assign n8298 = n8295 | n8297;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:842:89  */
  assign n8299 = exe_engine[23:19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:842:130  */
  assign n8301 = n8299 != 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:842:72  */
  assign n8302 = n8298 | n8301;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:842:9  */
  assign n8304 = n8302 ? 1'b1 : 1'b0;
  assign n8306 = {n8265, n8260, n8241, n8233, n8230, n8207, n8197, n8017, n8011, n7997, n7968};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8307 = 1'b0;
      11'b01000000000: n8307 = 1'b0;
      11'b00100000000: n8307 = 1'b0;
      11'b00010000000: n8307 = 1'b0;
      11'b00001000000: n8307 = n8225;
      11'b00000100000: n8307 = 1'b0;
      11'b00000010000: n8307 = 1'b0;
      11'b00000001000: n8307 = 1'b1;
      11'b00000000100: n8307 = 1'b0;
      11'b00000000010: n8307 = 1'b0;
      11'b00000000001: n8307 = 1'b0;
      default: n8307 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8308 = 1'b0;
      11'b01000000000: n8308 = 1'b0;
      11'b00100000000: n8308 = 1'b0;
      11'b00010000000: n8308 = 1'b0;
      11'b00001000000: n8308 = 1'b0;
      11'b00000100000: n8308 = 1'b0;
      11'b00000010000: n8308 = 1'b0;
      11'b00000001000: n8308 = 1'b0;
      11'b00000000100: n8308 = 1'b0;
      11'b00000000010: n8308 = 1'b0;
      11'b00000000001: n8308 = n7958;
      default: n8308 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8309 = n8263;
      11'b01000000000: n8309 = n8256;
      11'b00100000000: n8309 = 4'b1011;
      11'b00010000000: n8309 = 4'b0000;
      11'b00001000000: n8309 = n8226;
      11'b00000100000: n8309 = n8203;
      11'b00000010000: n8309 = n8178;
      11'b00000001000: n8309 = 4'b1000;
      11'b00000000100: n8309 = 4'b0011;
      11'b00000000010: n8309 = n7994;
      11'b00000000001: n8309 = n7961;
      default: n8309 = n8290;
    endcase
  assign n8310 = {n7852, n7851, n7850};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8311 = n8310;
      11'b01000000000: n8311 = n8310;
      11'b00100000000: n8311 = n8310;
      11'b00010000000: n8311 = n8310;
      11'b00001000000: n8311 = n8310;
      11'b00000100000: n8311 = n8310;
      11'b00000010000: n8311 = n8310;
      11'b00000001000: n8311 = n8310;
      11'b00000000100: n8311 = n8310;
      11'b00000000010: n8311 = n8310;
      11'b00000000001: n8311 = n7964;
      default: n8311 = n8310;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8312 = n7853;
      11'b01000000000: n8312 = n7853;
      11'b00100000000: n8312 = n7853;
      11'b00010000000: n8312 = n7853;
      11'b00001000000: n8312 = n8227;
      11'b00000100000: n8312 = n7853;
      11'b00000010000: n8312 = n8020;
      11'b00000001000: n8312 = n7853;
      11'b00000000100: n8312 = n8007;
      11'b00000000010: n8312 = n7990;
      11'b00000000001: n8312 = n7853;
      default: n8312 = n7853;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8313 = 32'b00000000000000000000000000000000;
      11'b01000000000: n8313 = 32'b00000000000000000000000000000000;
      11'b00100000000: n8313 = 32'b00000000000000000000000000000000;
      11'b00010000000: n8313 = 32'b00000000000000000000000000000000;
      11'b00001000000: n8313 = n8210;
      11'b00000100000: n8313 = 32'b00000000000000000000000000000000;
      11'b00000010000: n8313 = 32'b00000000000000000000000000000000;
      11'b00000001000: n8313 = 32'b00000000000000000000000000000000;
      11'b00000000100: n8313 = 32'b00000000000000000000000000000000;
      11'b00000000010: n8313 = 32'b00000000000000000000000000000000;
      11'b00000000001: n8313 = 32'b00000000000000000000000000000000;
      default: n8313 = 32'b00000000000000000000000000000000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8314 = 1'b0;
      11'b01000000000: n8314 = 1'b0;
      11'b00100000000: n8314 = 1'b0;
      11'b00010000000: n8314 = 1'b0;
      11'b00001000000: n8314 = 1'b0;
      11'b00000100000: n8314 = 1'b0;
      11'b00000010000: n8314 = 1'b0;
      11'b00000001000: n8314 = 1'b0;
      11'b00000000100: n8314 = 1'b0;
      11'b00000000010: n8314 = n7995;
      11'b00000000001: n8314 = 1'b0;
      default: n8314 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8315 = 1'b0;
      11'b01000000000: n8315 = 1'b0;
      11'b00100000000: n8315 = 1'b0;
      11'b00010000000: n8315 = 1'b0;
      11'b00001000000: n8315 = 1'b0;
      11'b00000100000: n8315 = 1'b0;
      11'b00000010000: n8315 = 1'b0;
      11'b00000001000: n8315 = 1'b0;
      11'b00000000100: n8315 = 1'b1;
      11'b00000000010: n8315 = 1'b0;
      11'b00000000001: n8315 = 1'b0;
      default: n8315 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8316 = 1'b0;
      11'b01000000000: n8316 = 1'b0;
      11'b00100000000: n8316 = 1'b0;
      11'b00010000000: n8316 = 1'b0;
      11'b00001000000: n8316 = 1'b0;
      11'b00000100000: n8316 = 1'b0;
      11'b00000010000: n8316 = pmp_fault_i;
      11'b00000001000: n8316 = 1'b0;
      11'b00000000100: n8316 = 1'b0;
      11'b00000000010: n8316 = 1'b0;
      11'b00000000001: n8316 = n7965;
      default: n8316 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8317 = 1'b0;
      11'b01000000000: n8317 = 1'b0;
      11'b00100000000: n8317 = 1'b0;
      11'b00010000000: n8317 = 1'b0;
      11'b00001000000: n8317 = n8228;
      11'b00000100000: n8317 = 1'b0;
      11'b00000010000: n8317 = 1'b0;
      11'b00000001000: n8317 = 1'b0;
      11'b00000000100: n8317 = 1'b0;
      11'b00000000010: n8317 = 1'b0;
      11'b00000000001: n8317 = 1'b0;
      default: n8317 = 1'b0;
    endcase
  assign n8318 = {1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8319 = n8318;
      11'b01000000000: n8319 = n8318;
      11'b00100000000: n8319 = n8318;
      11'b00010000000: n8319 = n8318;
      11'b00001000000: n8319 = n8318;
      11'b00000100000: n8319 = n8318;
      11'b00000010000: n8319 = n8318;
      11'b00000001000: n8319 = n8318;
      11'b00000000100: n8319 = n8318;
      11'b00000000010: n8319 = n8318;
      11'b00000000001: n8319 = n8318;
      default: n8319 = n8293;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8320 = 1'b0;
      11'b01000000000: n8320 = 1'b0;
      11'b00100000000: n8320 = 1'b0;
      11'b00010000000: n8320 = 1'b0;
      11'b00001000000: n8320 = 1'b0;
      11'b00000100000: n8320 = 1'b0;
      11'b00000010000: n8320 = 1'b0;
      11'b00000001000: n8320 = 1'b0;
      11'b00000000100: n8320 = 1'b0;
      11'b00000000010: n8320 = 1'b0;
      11'b00000000001: n8320 = n7966;
      default: n8320 = 1'b0;
    endcase
  assign n8321 = n7870[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8322 = n8321;
      11'b01000000000: n8322 = n8321;
      11'b00100000000: n8322 = n8321;
      11'b00010000000: n8322 = n8321;
      11'b00001000000: n8322 = n8321;
      11'b00000100000: n8322 = n8321;
      11'b00000010000: n8322 = n8180;
      11'b00000001000: n8322 = n8321;
      11'b00000000100: n8322 = n8321;
      11'b00000000010: n8322 = n8321;
      11'b00000000001: n8322 = n8321;
      default: n8322 = n8321;
    endcase
  assign n8323 = n7870[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8324 = n8323;
      11'b01000000000: n8324 = n8258;
      11'b00100000000: n8324 = n8323;
      11'b00010000000: n8324 = n8323;
      11'b00001000000: n8324 = n8211;
      11'b00000100000: n8324 = n8205;
      11'b00000010000: n8324 = n8182;
      11'b00000001000: n8324 = n8323;
      11'b00000000100: n8324 = n8323;
      11'b00000000010: n8324 = n8323;
      11'b00000000001: n8324 = n8323;
      default: n8324 = 1'b1;
    endcase
  assign n8325 = n7870[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8326 = n8325;
      11'b01000000000: n8326 = n8325;
      11'b00100000000: n8326 = n8325;
      11'b00010000000: n8326 = n8325;
      11'b00001000000: n8326 = n8325;
      11'b00000100000: n8326 = n8325;
      11'b00000010000: n8326 = n8325;
      11'b00000001000: n8326 = 1'b0;
      11'b00000000100: n8326 = n8325;
      11'b00000000010: n8326 = n8325;
      11'b00000000001: n8326 = n8325;
      default: n8326 = n8325;
    endcase
  assign n8327 = n7870[20:18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8328 = n8327;
      11'b01000000000: n8328 = n8327;
      11'b00100000000: n8328 = n8327;
      11'b00010000000: n8328 = n8327;
      11'b00001000000: n8328 = n8327;
      11'b00000100000: n8328 = 3'b010;
      11'b00000010000: n8328 = n8184;
      11'b00000001000: n8328 = n8327;
      11'b00000000100: n8328 = n8327;
      11'b00000000010: n8328 = n8327;
      11'b00000000001: n8328 = n8327;
      default: n8328 = n8327;
    endcase
  assign n8329 = n7870[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8330 = n8329;
      11'b01000000000: n8330 = n8329;
      11'b00100000000: n8330 = n8329;
      11'b00010000000: n8330 = n8329;
      11'b00001000000: n8330 = n8329;
      11'b00000100000: n8330 = n8329;
      11'b00000010000: n8330 = n8186;
      11'b00000001000: n8330 = n8329;
      11'b00000000100: n8330 = n8329;
      11'b00000000010: n8330 = n8329;
      11'b00000000001: n8330 = n8329;
      default: n8330 = n8329;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8331 = n7883;
      11'b01000000000: n8331 = n7883;
      11'b00100000000: n8331 = n7883;
      11'b00010000000: n8331 = n7883;
      11'b00001000000: n8331 = n7883;
      11'b00000100000: n8331 = n7883;
      11'b00000010000: n8331 = n7883;
      11'b00000001000: n8331 = n7883;
      11'b00000000100: n8331 = n7883;
      11'b00000000010: n8331 = n7883;
      11'b00000000001: n8331 = 1'b1;
      default: n8331 = n7883;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8332 = n7914;
      11'b01000000000: n8332 = n7914;
      11'b00100000000: n8332 = n7914;
      11'b00010000000: n8332 = n7914;
      11'b00001000000: n8332 = n7914;
      11'b00000100000: n8332 = n7914;
      11'b00000010000: n8332 = n7914;
      11'b00000001000: n8332 = n7914;
      11'b00000000100: n8332 = n7914;
      11'b00000000010: n8332 = n7914;
      11'b00000000001: n8332 = 1'b1;
      default: n8332 = n7914;
    endcase
  assign n8333 = n7870[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8334 = n8333;
      11'b01000000000: n8334 = n8333;
      11'b00100000000: n8334 = n8333;
      11'b00010000000: n8334 = n8333;
      11'b00001000000: n8334 = n8333;
      11'b00000100000: n8334 = n8333;
      11'b00000010000: n8334 = n8188;
      11'b00000001000: n8334 = n8333;
      11'b00000000100: n8334 = n8333;
      11'b00000000010: n8334 = n8333;
      11'b00000000001: n8334 = n8333;
      default: n8334 = n8333;
    endcase
  assign n8335 = n7870[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8336 = n8335;
      11'b01000000000: n8336 = n8335;
      11'b00100000000: n8336 = n8335;
      11'b00010000000: n8336 = n8335;
      11'b00001000000: n8336 = n8335;
      11'b00000100000: n8336 = n8335;
      11'b00000010000: n8336 = n8190;
      11'b00000001000: n8336 = n8335;
      11'b00000000100: n8336 = n8335;
      11'b00000000010: n8336 = n8335;
      11'b00000000001: n8336 = n8335;
      default: n8336 = n8335;
    endcase
  assign n8337 = n7870[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8338 = n8337;
      11'b01000000000: n8338 = n8337;
      11'b00100000000: n8338 = n8337;
      11'b00010000000: n8338 = n8337;
      11'b00001000000: n8338 = n8337;
      11'b00000100000: n8338 = n8337;
      11'b00000010000: n8338 = n8192;
      11'b00000001000: n8338 = n8337;
      11'b00000000100: n8338 = n8337;
      11'b00000000010: n8338 = n8337;
      11'b00000000001: n8338 = n8337;
      default: n8338 = n8337;
    endcase
  assign n8339 = n7870[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8340 = n8339;
      11'b01000000000: n8340 = n8339;
      11'b00100000000: n8340 = n8238;
      11'b00010000000: n8340 = n8339;
      11'b00001000000: n8340 = n8339;
      11'b00000100000: n8340 = n8339;
      11'b00000010000: n8340 = n8339;
      11'b00000001000: n8340 = n8339;
      11'b00000000100: n8340 = n8339;
      11'b00000000010: n8340 = n8339;
      11'b00000000001: n8340 = n8339;
      default: n8340 = n8339;
    endcase
  assign n8341 = n7870[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8342 = n8341;
      11'b01000000000: n8342 = n8341;
      11'b00100000000: n8342 = n8341;
      11'b00010000000: n8342 = n8341;
      11'b00001000000: n8342 = n8341;
      11'b00000100000: n8342 = n8341;
      11'b00000010000: n8342 = n8194;
      11'b00000001000: n8342 = n8341;
      11'b00000000100: n8342 = n8341;
      11'b00000000010: n8342 = n8341;
      11'b00000000001: n8342 = n8341;
      default: n8342 = n8341;
    endcase
  assign n8346 = n7870[16:2]; // extract
  assign n8351 = n7870[58:32]; // extract
  assign n8352 = n7870[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8353 = 1'b0;
      11'b01000000000: n8353 = 1'b0;
      11'b00100000000: n8353 = 1'b0;
      11'b00010000000: n8353 = 1'b0;
      11'b00001000000: n8353 = 1'b0;
      11'b00000100000: n8353 = 1'b0;
      11'b00000010000: n8353 = 1'b0;
      11'b00000001000: n8353 = 1'b0;
      11'b00000000100: n8353 = 1'b0;
      11'b00000000010: n8353 = 1'b0;
      11'b00000000001: n8353 = 1'b0;
      default: n8353 = n8304;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:636:5  */
  always @*
    case (n8306)
      11'b10000000000: n8354 = 1'b0;
      11'b01000000000: n8354 = 1'b0;
      11'b00100000000: n8354 = 1'b0;
      11'b00010000000: n8354 = 1'b0;
      11'b00001000000: n8354 = 1'b0;
      11'b00000100000: n8354 = 1'b0;
      11'b00000010000: n8354 = n8195;
      11'b00000001000: n8354 = 1'b0;
      11'b00000000100: n8354 = 1'b0;
      11'b00000000010: n8354 = 1'b0;
      11'b00000000001: n8354 = 1'b0;
      default: n8354 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:856:31  */
  assign n8356 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:858:31  */
  assign n8357 = ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:858:59  */
  assign n8358 = trap_ctrl[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:858:45  */
  assign n8359 = ~n8358;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:858:40  */
  assign n8360 = n8357 & n8359;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:859:39  */
  assign n8361 = exe_engine[23:19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:860:39  */
  assign n8362 = exe_engine[28:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:861:39  */
  assign n8363 = exe_engine[15:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:862:31  */
  assign n8364 = ctrl[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:864:31  */
  assign n8365 = ctrl[20:18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:865:31  */
  assign n8366 = ctrl[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:866:31  */
  assign n8367 = ctrl[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:867:31  */
  assign n8368 = ctrl[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:868:31  */
  assign n8369 = ctrl[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:869:31  */
  assign n8370 = ctrl[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:870:31  */
  assign n8371 = ctrl[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:871:31  */
  assign n8372 = ctrl[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:873:31  */
  assign n8373 = ctrl[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:874:31  */
  assign n8374 = ctrl[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:875:47  */
  assign n8376 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:875:53  */
  assign n8378 = n8376 == 4'b1010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:875:30  */
  assign n8379 = n8378 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:876:31  */
  assign n8381 = ctrl[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:877:30  */
  assign n8382 = csr[114]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:877:52  */
  assign n8383 = csr[115]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:877:42  */
  assign n8384 = n8383 ? n8382 : n8385;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:877:81  */
  assign n8385 = csr[137]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:879:39  */
  assign n8386 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:880:39  */
  assign n8387 = exe_engine[35:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:883:30  */
  assign n8388 = csr[137]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:885:36  */
  assign n8389 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:886:37  */
  assign n8390 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:897:16  */
  assign n8392 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:900:22  */
  assign n8394 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:900:28  */
  assign n8396 = n8394 == 4'b0110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:901:64  */
  assign n8398 = monitor_cnt + 10'b0000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:900:7  */
  assign n8400 = n8396 ? n8398 : 10'b0000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:909:29  */
  assign n8405 = monitor_cnt[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:918:32  */
  assign n8408 = exe_engine[35:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:926:7  */
  assign n8412 = n8408 == 12'b100000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:926:26  */
  assign n8414 = n8408 == 12'b100000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:926:26  */
  assign n8415 = n8412 | n8414;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:926:42  */
  assign n8417 = n8408 == 12'b100000000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:926:42  */
  assign n8418 = n8415 | n8417;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:926:58  */
  assign n8420 = n8408 == 12'b100000000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:926:58  */
  assign n8421 = n8418 | n8420;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:930:7  */
  assign n8425 = n8408 == 12'b000000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:930:25  */
  assign n8427 = n8408 == 12'b000000000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:930:25  */
  assign n8428 = n8425 | n8427;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:930:37  */
  assign n8430 = n8408 == 12'b000000000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:930:37  */
  assign n8431 = n8428 | n8430;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:7  */
  assign n8434 = n8408 == 12'b001100000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:28  */
  assign n8436 = n8408 == 12'b001100010000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:28  */
  assign n8437 = n8434 | n8436;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:50  */
  assign n8439 = n8408 == 12'b001100000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:50  */
  assign n8440 = n8437 | n8439;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:68  */
  assign n8442 = n8408 == 12'b001100000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:68  */
  assign n8443 = n8440 | n8442;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:86  */
  assign n8445 = n8408 == 12'b001100000101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:86  */
  assign n8446 = n8443 | n8445;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:101  */
  assign n8448 = n8408 == 12'b001101000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:934:101  */
  assign n8449 = n8446 | n8448;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:28  */
  assign n8451 = n8408 == 12'b001101000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:28  */
  assign n8452 = n8449 | n8451;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:50  */
  assign n8454 = n8408 == 12'b001101000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:50  */
  assign n8455 = n8452 | n8454;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:68  */
  assign n8457 = n8408 == 12'b001101000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:68  */
  assign n8458 = n8455 | n8457;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:86  */
  assign n8460 = n8408 == 12'b001101000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:86  */
  assign n8461 = n8458 | n8460;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:101  */
  assign n8463 = n8408 == 12'b001101001010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:935:101  */
  assign n8464 = n8461 | n8463;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:28  */
  assign n8466 = n8408 == 12'b001100100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:28  */
  assign n8467 = n8464 | n8466;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:50  */
  assign n8469 = n8408 == 12'b111100010001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:50  */
  assign n8470 = n8467 | n8469;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:68  */
  assign n8472 = n8408 == 12'b111100010010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:68  */
  assign n8473 = n8470 | n8472;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:86  */
  assign n8475 = n8408 == 12'b111100010011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:86  */
  assign n8476 = n8473 | n8475;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:101  */
  assign n8478 = n8408 == 12'b111100010100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:936:101  */
  assign n8479 = n8476 | n8478;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:937:28  */
  assign n8481 = n8408 == 12'b111100010101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:937:28  */
  assign n8482 = n8479 | n8481;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:937:50  */
  assign n8484 = n8408 == 12'b111111000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:937:50  */
  assign n8485 = n8482 | n8484;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:937:68  */
  assign n8487 = n8408 == 12'b101111000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:937:68  */
  assign n8488 = n8485 | n8487;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:937:86  */
  assign n8490 = n8408 == 12'b101111000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:937:86  */
  assign n8491 = n8488 | n8490;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:941:7  */
  assign n8495 = n8408 == 12'b001100000110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:941:29  */
  assign n8497 = n8408 == 12'b001100001010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:941:29  */
  assign n8498 = n8495 | n8497;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:941:45  */
  assign n8500 = n8408 == 12'b001100011010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:941:45  */
  assign n8501 = n8498 | n8500;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:7  */
  assign n8505 = n8408 == 12'b001110100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:28  */
  assign n8507 = n8408 == 12'b001110100001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:28  */
  assign n8508 = n8505 | n8507;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:46  */
  assign n8510 = n8408 == 12'b001110100010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:46  */
  assign n8511 = n8508 | n8510;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:64  */
  assign n8513 = n8408 == 12'b001110100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:64  */
  assign n8514 = n8511 | n8513;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:82  */
  assign n8516 = n8408 == 12'b001110110000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:945:82  */
  assign n8517 = n8514 | n8516;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:946:28  */
  assign n8519 = n8408 == 12'b001110110001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:946:28  */
  assign n8520 = n8517 | n8519;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:946:46  */
  assign n8522 = n8408 == 12'b001110110010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:946:46  */
  assign n8523 = n8520 | n8522;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:946:64  */
  assign n8525 = n8408 == 12'b001110110011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:946:64  */
  assign n8526 = n8523 | n8525;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:946:82  */
  assign n8528 = n8408 == 12'b001110110100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:946:82  */
  assign n8529 = n8526 | n8528;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:947:28  */
  assign n8531 = n8408 == 12'b001110110101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:947:28  */
  assign n8532 = n8529 | n8531;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:947:46  */
  assign n8534 = n8408 == 12'b001110110110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:947:46  */
  assign n8535 = n8532 | n8534;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:947:64  */
  assign n8537 = n8408 == 12'b001110110111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:947:64  */
  assign n8538 = n8535 | n8537;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:947:82  */
  assign n8540 = n8408 == 12'b001110111000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:947:82  */
  assign n8541 = n8538 | n8540;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:948:28  */
  assign n8543 = n8408 == 12'b001110111001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:948:28  */
  assign n8544 = n8541 | n8543;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:948:46  */
  assign n8546 = n8408 == 12'b001110111010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:948:46  */
  assign n8547 = n8544 | n8546;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:948:64  */
  assign n8549 = n8408 == 12'b001110111011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:948:64  */
  assign n8550 = n8547 | n8549;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:948:82  */
  assign n8552 = n8408 == 12'b001110111100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:948:82  */
  assign n8553 = n8550 | n8552;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:949:28  */
  assign n8555 = n8408 == 12'b001110111101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:949:28  */
  assign n8556 = n8553 | n8555;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:949:46  */
  assign n8558 = n8408 == 12'b001110111110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:949:46  */
  assign n8559 = n8556 | n8558;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:949:64  */
  assign n8561 = n8408 == 12'b001110111111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:949:64  */
  assign n8562 = n8559 | n8561;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:7  */
  assign n8566 = n8408 == 12'b101100000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:33  */
  assign n8568 = n8408 == 12'b101100000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:33  */
  assign n8569 = n8566 | n8568;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:56  */
  assign n8571 = n8408 == 12'b101100000101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:56  */
  assign n8572 = n8569 | n8571;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:79  */
  assign n8574 = n8408 == 12'b101100000110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:79  */
  assign n8575 = n8572 | n8574;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:102  */
  assign n8577 = n8408 == 12'b101100000111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:102  */
  assign n8578 = n8575 | n8577;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:125  */
  assign n8580 = n8408 == 12'b101100001000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:953:125  */
  assign n8581 = n8578 | n8580;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:33  */
  assign n8583 = n8408 == 12'b101100001001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:33  */
  assign n8584 = n8581 | n8583;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:56  */
  assign n8586 = n8408 == 12'b101100001010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:56  */
  assign n8587 = n8584 | n8586;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:79  */
  assign n8589 = n8408 == 12'b101100001011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:79  */
  assign n8590 = n8587 | n8589;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:102  */
  assign n8592 = n8408 == 12'b101100001100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:102  */
  assign n8593 = n8590 | n8592;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:125  */
  assign n8595 = n8408 == 12'b101100001101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:954:125  */
  assign n8596 = n8593 | n8595;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:955:33  */
  assign n8598 = n8408 == 12'b101100001110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:955:33  */
  assign n8599 = n8596 | n8598;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:955:56  */
  assign n8601 = n8408 == 12'b101100001111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:955:56  */
  assign n8602 = n8599 | n8601;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:955:79  */
  assign n8604 = n8408 == 12'b101110000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:955:79  */
  assign n8605 = n8602 | n8604;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:33  */
  assign n8607 = n8408 == 12'b101110000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:33  */
  assign n8608 = n8605 | n8607;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:56  */
  assign n8610 = n8408 == 12'b101110000101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:56  */
  assign n8611 = n8608 | n8610;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:79  */
  assign n8613 = n8408 == 12'b101110000110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:79  */
  assign n8614 = n8611 | n8613;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:102  */
  assign n8616 = n8408 == 12'b101110000111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:102  */
  assign n8617 = n8614 | n8616;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:125  */
  assign n8619 = n8408 == 12'b101110001000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:956:125  */
  assign n8620 = n8617 | n8619;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:33  */
  assign n8622 = n8408 == 12'b101110001001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:33  */
  assign n8623 = n8620 | n8622;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:56  */
  assign n8625 = n8408 == 12'b101110001010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:56  */
  assign n8626 = n8623 | n8625;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:79  */
  assign n8628 = n8408 == 12'b101110001011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:79  */
  assign n8629 = n8626 | n8628;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:102  */
  assign n8631 = n8408 == 12'b101110001100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:102  */
  assign n8632 = n8629 | n8631;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:125  */
  assign n8634 = n8408 == 12'b101110001101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:957:125  */
  assign n8635 = n8632 | n8634;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:958:33  */
  assign n8637 = n8408 == 12'b101110001110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:958:33  */
  assign n8638 = n8635 | n8637;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:958:56  */
  assign n8640 = n8408 == 12'b101110001111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:958:56  */
  assign n8641 = n8638 | n8640;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:958:79  */
  assign n8643 = n8408 == 12'b001100100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:958:79  */
  assign n8644 = n8641 | n8643;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:33  */
  assign n8646 = n8408 == 12'b001100100100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:33  */
  assign n8647 = n8644 | n8646;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:56  */
  assign n8649 = n8408 == 12'b001100100101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:56  */
  assign n8650 = n8647 | n8649;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:79  */
  assign n8652 = n8408 == 12'b001100100110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:79  */
  assign n8653 = n8650 | n8652;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:102  */
  assign n8655 = n8408 == 12'b001100100111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:102  */
  assign n8656 = n8653 | n8655;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:125  */
  assign n8658 = n8408 == 12'b001100101000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:959:125  */
  assign n8659 = n8656 | n8658;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:33  */
  assign n8661 = n8408 == 12'b001100101001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:33  */
  assign n8662 = n8659 | n8661;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:56  */
  assign n8664 = n8408 == 12'b001100101010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:56  */
  assign n8665 = n8662 | n8664;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:79  */
  assign n8667 = n8408 == 12'b001100101011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:79  */
  assign n8668 = n8665 | n8667;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:102  */
  assign n8670 = n8408 == 12'b001100101100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:102  */
  assign n8671 = n8668 | n8670;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:125  */
  assign n8673 = n8408 == 12'b001100101101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:960:125  */
  assign n8674 = n8671 | n8673;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:961:33  */
  assign n8676 = n8408 == 12'b001100101110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:961:33  */
  assign n8677 = n8674 | n8676;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:961:56  */
  assign n8679 = n8408 == 12'b001100101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:961:56  */
  assign n8680 = n8677 | n8679;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:7  */
  assign n8684 = n8408 == 12'b110000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:24  */
  assign n8686 = n8408 == 12'b101100000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:24  */
  assign n8687 = n8684 | n8686;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:39  */
  assign n8689 = n8408 == 12'b110000000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:39  */
  assign n8690 = n8687 | n8689;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:55  */
  assign n8692 = n8408 == 12'b101100000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:55  */
  assign n8693 = n8690 | n8692;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:72  */
  assign n8695 = n8408 == 12'b110010000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:72  */
  assign n8696 = n8693 | n8695;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:87  */
  assign n8698 = n8408 == 12'b101110000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:87  */
  assign n8699 = n8696 | n8698;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:103  */
  assign n8701 = n8408 == 12'b110010000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:103  */
  assign n8702 = n8699 | n8701;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:120  */
  assign n8704 = n8408 == 12'b101110000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:965:120  */
  assign n8705 = n8702 | n8704;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:969:7  */
  assign n8709 = n8408 == 12'b011110110000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:969:23  */
  assign n8711 = n8408 == 12'b011110110001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:969:23  */
  assign n8712 = n8709 | n8711;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:969:35  */
  assign n8714 = n8408 == 12'b011110110010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:969:35  */
  assign n8715 = n8712 | n8714;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:973:7  */
  assign n8719 = n8408 == 12'b011110100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:973:26  */
  assign n8721 = n8408 == 12'b011110100001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:973:26  */
  assign n8722 = n8719 | n8721;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:973:41  */
  assign n8724 = n8408 == 12'b011110100010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:973:41  */
  assign n8725 = n8722 | n8724;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:973:56  */
  assign n8727 = n8408 == 12'b011110100100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:973:56  */
  assign n8728 = n8725 | n8727;
  assign n8730 = {n8728, n8715, n8705, n8680, n8562, n8501, n8491, n8431, n8421};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:923:5  */
  always @*
    case (n8730)
      9'b100000000: n8731 = 1'b1;
      9'b010000000: n8731 = 1'b1;
      9'b001000000: n8731 = 1'b1;
      9'b000100000: n8731 = 1'b0;
      9'b000010000: n8731 = 1'b0;
      9'b000001000: n8731 = 1'b1;
      9'b000000100: n8731 = 1'b1;
      9'b000000010: n8731 = 1'b0;
      9'b000000001: n8731 = 1'b0;
      default: n8731 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:985:19  */
  assign n8732 = exe_engine[35:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:985:34  */
  assign n8734 = n8732 == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:986:23  */
  assign n8735 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:986:70  */
  assign n8737 = n8735 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:987:23  */
  assign n8738 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:987:70  */
  assign n8740 = n8738 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:986:89  */
  assign n8741 = n8737 | n8740;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:988:23  */
  assign n8742 = exe_engine[23:19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:988:64  */
  assign n8744 = n8742 != 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:987:89  */
  assign n8745 = n8741 | n8744;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:985:42  */
  assign n8746 = n8745 & n8734;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:985:5  */
  assign n8749 = n8746 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:997:19  */
  assign n8750 = exe_engine[35:28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:997:33  */
  assign n8752 = n8750 == 8'b01111011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:997:60  */
  assign n8754 = 1'b1 & n8752;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:998:40  */
  assign n8755 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:998:44  */
  assign n8756 = ~n8755;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:998:24  */
  assign n8757 = n8756 & n8754;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1000:53  */
  assign n8759 = csr[137]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1000:67  */
  assign n8760 = ~n8759;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1000:44  */
  assign n8762 = n8760 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1001:22  */
  assign n8763 = exe_engine[35:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1001:36  */
  assign n8765 = n8763 == 4'b1100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1000:74  */
  assign n8766 = n8765 & n8762;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1002:24  */
  assign n8767 = exe_engine[25:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1002:37  */
  assign n8769 = n8767 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1002:73  */
  assign n8770 = csr[304]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1002:87  */
  assign n8771 = ~n8770;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1002:64  */
  assign n8772 = n8771 & n8769;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1003:24  */
  assign n8773 = exe_engine[25:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1003:37  */
  assign n8775 = n8773 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1003:75  */
  assign n8776 = csr[305]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1003:89  */
  assign n8777 = ~n8776;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1003:66  */
  assign n8778 = n8777 & n8775;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1002:95  */
  assign n8779 = n8772 | n8778;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1001:64  */
  assign n8780 = n8779 & n8766;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1005:22  */
  assign n8782 = exe_engine[33:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1005:35  */
  assign n8784 = n8782 != 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1005:53  */
  assign n8785 = csr[137]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1005:67  */
  assign n8786 = ~n8785;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1005:44  */
  assign n8787 = n8786 & n8784;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1005:5  */
  assign n8790 = n8787 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1000:5  */
  assign n8791 = n8780 ? 1'b0 : n8790;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:997:5  */
  assign n8792 = n8757 ? 1'b0 : n8791;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1019:23  */
  assign n8795 = exe_engine[10:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1021:7  */
  assign n8797 = n8795 == 7'b0110111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1021:25  */
  assign n8799 = n8795 == 7'b0010111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1021:25  */
  assign n8800 = n8797 | n8799;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1021:42  */
  assign n8802 = n8795 == 7'b1101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1021:42  */
  assign n8803 = n8800 | n8802;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1025:26  */
  assign n8804 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1025:73  */
  assign n8806 = n8804 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1025:9  */
  assign n8809 = n8806 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1024:7  */
  assign n8811 = n8795 == 7'b1100111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1030:27  */
  assign n8812 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:11  */
  assign n8814 = n8812 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:29  */
  assign n8816 = n8812 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:29  */
  assign n8817 = n8814 | n8816;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:44  */
  assign n8819 = n8812 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:44  */
  assign n8820 = n8817 | n8819;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:59  */
  assign n8822 = n8812 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:59  */
  assign n8823 = n8820 | n8822;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:74  */
  assign n8825 = n8812 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:74  */
  assign n8826 = n8823 | n8825;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:90  */
  assign n8828 = n8812 == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1031:90  */
  assign n8829 = n8826 | n8828;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1030:9  */
  always @*
    case (n8829)
      1'b1: n8832 = 1'b0;
      default: n8832 = 1'b1;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1029:7  */
  assign n8834 = n8795 == 7'b1100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1036:27  */
  assign n8835 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:11  */
  assign n8837 = n8835 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:28  */
  assign n8839 = n8835 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:28  */
  assign n8840 = n8837 | n8839;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:42  */
  assign n8842 = n8835 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:42  */
  assign n8843 = n8840 | n8842;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:56  */
  assign n8845 = n8835 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:56  */
  assign n8846 = n8843 | n8845;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:71  */
  assign n8848 = n8835 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1037:71  */
  assign n8849 = n8846 | n8848;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1036:9  */
  always @*
    case (n8849)
      1'b1: n8852 = 1'b0;
      default: n8852 = 1'b1;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1035:7  */
  assign n8854 = n8795 == 7'b0000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1042:27  */
  assign n8855 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1043:11  */
  assign n8857 = n8855 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1043:28  */
  assign n8859 = n8855 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1043:28  */
  assign n8860 = n8857 | n8859;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1043:42  */
  assign n8862 = n8855 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1043:42  */
  assign n8863 = n8860 | n8862;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1042:9  */
  always @*
    case (n8863)
      1'b1: n8866 = 1'b0;
      default: n8866 = 1'b1;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1041:7  */
  assign n8868 = n8795 == 7'b0100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1047:7  */
  assign n8870 = n8795 == 7'b0101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:7  */
  assign n8872 = n8795 == 7'b0110011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:25  */
  assign n8874 = n8795 == 7'b0010011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:25  */
  assign n8875 = n8872 | n8874;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:41  */
  assign n8877 = n8795 == 7'b1010011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:41  */
  assign n8878 = n8875 | n8877;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:56  */
  assign n8880 = n8795 == 7'b0001011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:56  */
  assign n8881 = n8878 | n8880;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:73  */
  assign n8883 = n8795 == 7'b0101011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1055:73  */
  assign n8884 = n8881 | n8883;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1059:26  */
  assign n8885 = exe_engine[18:17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1059:75  */
  assign n8887 = n8885 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1059:9  */
  assign n8890 = n8887 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1058:7  */
  assign n8892 = n8795 == 7'b0001111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1064:26  */
  assign n8893 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1064:73  */
  assign n8895 = n8893 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1065:28  */
  assign n8896 = exe_engine[23:19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1065:69  */
  assign n8898 = n8896 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1065:98  */
  assign n8899 = exe_engine[15:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1065:137  */
  assign n8901 = n8899 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1065:80  */
  assign n8902 = n8901 & n8898;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1066:31  */
  assign n8903 = exe_engine[35:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1067:15  */
  assign n8905 = n8903 == 12'b000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1068:15  */
  assign n8907 = n8903 == 12'b000000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1069:64  */
  assign n8908 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1069:56  */
  assign n8909 = ~n8908;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1069:89  */
  assign n8910 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1069:75  */
  assign n8911 = n8909 | n8910;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1069:15  */
  assign n8913 = n8903 == 12'b001100000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1070:70  */
  assign n8914 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1070:55  */
  assign n8915 = ~n8914;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1070:15  */
  assign n8917 = n8903 == 12'b011110110010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1071:64  */
  assign n8918 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1071:56  */
  assign n8919 = ~n8918;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1071:83  */
  assign n8920 = csr[116]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1071:75  */
  assign n8921 = n8919 & n8920;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1071:15  */
  assign n8923 = n8903 == 12'b000100000101;
  assign n8924 = {n8923, n8917, n8913, n8907, n8905};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1066:13  */
  always @*
    case (n8924)
      5'b10000: n8928 = n8921;
      5'b01000: n8928 = n8915;
      5'b00100: n8928 = n8911;
      5'b00010: n8928 = 1'b0;
      5'b00001: n8928 = 1'b0;
      default: n8928 = 1'b1;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1065:11  */
  assign n8930 = n8902 ? n8928 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1075:26  */
  assign n8932 = csr_valid == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1075:53  */
  assign n8933 = exe_engine[18:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1075:100  */
  assign n8935 = n8933 != 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1075:35  */
  assign n8936 = n8935 & n8932;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1075:9  */
  assign n8939 = n8936 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1064:9  */
  assign n8940 = n8895 ? n8930 : n8939;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1063:7  */
  assign n8942 = n8795 == 7'b1110011;
  assign n8943 = {n8942, n8892, n8884, n8870, n8868, n8854, n8834, n8811, n8803};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1019:5  */
  always @*
    case (n8943)
      9'b100000000: n8948 = n8940;
      9'b010000000: n8948 = n8890;
      9'b001000000: n8948 = 1'b0;
      9'b000100000: n8948 = 1'b1;
      9'b000010000: n8948 = n8866;
      9'b000001000: n8948 = n8852;
      9'b000000100: n8948 = n8832;
      9'b000000010: n8948 = n8809;
      9'b000000001: n8948 = 1'b0;
      default: n8948 = 1'b1;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1088:47  */
  assign n8952 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1088:53  */
  assign n8954 = n8952 == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1088:82  */
  assign n8955 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1088:88  */
  assign n8957 = n8955 == 4'b0110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1088:67  */
  assign n8958 = n8954 | n8957;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1089:55  */
  assign n8959 = monitor_exc | illegal_cmd;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1088:104  */
  assign n8960 = n8959 & n8958;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1088:29  */
  assign n8961 = n8960 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1100:16  */
  assign n8964 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1112:60  */
  assign n8967 = trap_ctrl[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1112:87  */
  assign n8968 = lsu_err_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1112:75  */
  assign n8969 = n8967 | n8968;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1112:117  */
  assign n8970 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1112:103  */
  assign n8971 = ~n8970;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1112:98  */
  assign n8972 = n8969 & n8971;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1113:60  */
  assign n8973 = trap_ctrl[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1113:87  */
  assign n8974 = lsu_err_i[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1113:75  */
  assign n8975 = n8973 | n8974;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1113:117  */
  assign n8976 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1113:103  */
  assign n8977 = ~n8976;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1113:98  */
  assign n8978 = n8975 & n8977;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1114:60  */
  assign n8979 = trap_ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1114:88  */
  assign n8980 = trap_ctrl[102]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1114:75  */
  assign n8981 = n8979 | n8980;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1114:117  */
  assign n8982 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1114:103  */
  assign n8983 = ~n8982;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1114:98  */
  assign n8984 = n8981 & n8983;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1117:61  */
  assign n8985 = trap_ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1117:89  */
  assign n8986 = lsu_err_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1117:77  */
  assign n8987 = n8985 | n8986;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1117:119  */
  assign n8988 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1117:105  */
  assign n8989 = ~n8988;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1117:100  */
  assign n8990 = n8987 & n8989;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1118:61  */
  assign n8991 = trap_ctrl[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1118:89  */
  assign n8992 = lsu_err_i[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1118:77  */
  assign n8993 = n8991 | n8992;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1118:119  */
  assign n8994 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1118:105  */
  assign n8995 = ~n8994;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1118:100  */
  assign n8996 = n8993 & n8995;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1119:61  */
  assign n8997 = trap_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1119:90  */
  assign n8998 = trap_ctrl[101]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1119:77  */
  assign n8999 = n8997 | n8998;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1119:119  */
  assign n9000 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1119:105  */
  assign n9001 = ~n9000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1119:100  */
  assign n9002 = n8999 & n9001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1122:61  */
  assign n9003 = trap_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1122:90  */
  assign n9004 = trap_ctrl[104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1122:77  */
  assign n9005 = n9003 | n9004;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1122:119  */
  assign n9006 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1122:105  */
  assign n9007 = ~n9006;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1122:100  */
  assign n9008 = n9005 & n9007;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1123:61  */
  assign n9009 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1123:90  */
  assign n9010 = trap_ctrl[103]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1123:77  */
  assign n9011 = n9009 | n9010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1123:119  */
  assign n9012 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1123:105  */
  assign n9013 = ~n9012;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1123:100  */
  assign n9014 = n9011 & n9013;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1127:59  */
  assign n9015 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1127:45  */
  assign n9016 = ~n9015;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1127:92  */
  assign n9017 = trap_ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1128:22  */
  assign n9018 = trap_ctrl[106]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1128:42  */
  assign n9019 = csr[426]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1128:34  */
  assign n9020 = ~n9019;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1128:29  */
  assign n9021 = n9018 & n9020;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1127:107  */
  assign n9022 = n9017 | n9021;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:22  */
  assign n9023 = trap_ctrl[105]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:42  */
  assign n9024 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:29  */
  assign n9025 = n9023 & n9024;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:66  */
  assign n9026 = csr[322]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:58  */
  assign n9027 = ~n9026;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:53  */
  assign n9028 = n9025 & n9027;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:100  */
  assign n9029 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:85  */
  assign n9030 = ~n9029;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:80  */
  assign n9031 = n9028 & n9030;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1128:58  */
  assign n9032 = n9022 | n9031;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:22  */
  assign n9033 = trap_ctrl[105]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:42  */
  assign n9034 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:34  */
  assign n9035 = ~n9034;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:29  */
  assign n9036 = n9033 & n9035;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:66  */
  assign n9037 = csr[323]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:58  */
  assign n9038 = ~n9037;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:53  */
  assign n9039 = n9036 & n9038;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:100  */
  assign n9040 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:85  */
  assign n9041 = ~n9040;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1130:80  */
  assign n9042 = n9039 & n9041;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1129:106  */
  assign n9043 = n9032 | n9042;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1127:70  */
  assign n9044 = n9016 & n9043;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1136:62  */
  assign n9045 = trap_ctrl[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1136:93  */
  assign n9046 = debug_ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1136:79  */
  assign n9047 = n9045 | n9046;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1136:124  */
  assign n9048 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1136:110  */
  assign n9049 = ~n9048;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1136:105  */
  assign n9050 = n9047 & n9049;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1137:62  */
  assign n9051 = trap_ctrl[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1137:93  */
  assign n9052 = debug_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1137:79  */
  assign n9053 = n9051 | n9052;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1137:124  */
  assign n9054 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1137:110  */
  assign n9055 = ~n9054;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1137:105  */
  assign n9056 = n9053 & n9055;
  assign n9057 = {n9056, n9050, n8990, n8996, n8972, n8978, n9044, n9008, n8984, n9014, n9002};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1146:16  */
  assign n9063 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1157:56  */
  assign n9067 = irq_machine_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1158:56  */
  assign n9068 = irq_machine_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1159:56  */
  assign n9069 = irq_machine_i[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1175:61  */
  assign n9072 = trap_ctrl[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1175:85  */
  assign n9073 = csr[117]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1175:77  */
  assign n9074 = n9072 & n9073;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1175:108  */
  assign n9075 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1175:141  */
  assign n9076 = trap_ctrl[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1175:120  */
  assign n9077 = n9075 & n9076;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1175:94  */
  assign n9078 = n9074 | n9077;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1176:61  */
  assign n9079 = trap_ctrl[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1176:85  */
  assign n9080 = csr[118]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1176:77  */
  assign n9081 = n9079 & n9080;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1176:108  */
  assign n9082 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1176:141  */
  assign n9083 = trap_ctrl[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1176:120  */
  assign n9084 = n9082 & n9083;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1176:94  */
  assign n9085 = n9081 | n9084;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1177:61  */
  assign n9086 = trap_ctrl[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1177:85  */
  assign n9087 = csr[119]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1177:77  */
  assign n9088 = n9086 & n9087;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1177:108  */
  assign n9089 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1177:141  */
  assign n9090 = trap_ctrl[34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1177:120  */
  assign n9091 = n9089 & n9090;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1177:94  */
  assign n9092 = n9088 | n9091;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9093 = trap_ctrl[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9094 = csr[120]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9095 = n9093 & n9094;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9096 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9097 = trap_ctrl[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9098 = n9096 & n9097;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9099 = n9095 | n9098;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9100 = trap_ctrl[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9101 = csr[121]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9102 = n9100 & n9101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9103 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9104 = trap_ctrl[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9105 = n9103 & n9104;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9106 = n9102 | n9105;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9107 = trap_ctrl[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9108 = csr[122]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9109 = n9107 & n9108;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9110 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9111 = trap_ctrl[38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9112 = n9110 & n9111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9113 = n9109 | n9112;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9114 = trap_ctrl[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9115 = csr[123]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9116 = n9114 & n9115;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9117 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9118 = trap_ctrl[39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9119 = n9117 & n9118;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9120 = n9116 | n9119;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9121 = trap_ctrl[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9122 = csr[124]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9123 = n9121 & n9122;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9124 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9125 = trap_ctrl[40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9126 = n9124 & n9125;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9127 = n9123 | n9126;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9128 = trap_ctrl[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9129 = csr[125]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9130 = n9128 & n9129;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9131 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9132 = trap_ctrl[41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9133 = n9131 & n9132;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9134 = n9130 | n9133;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9135 = trap_ctrl[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9136 = csr[126]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9137 = n9135 & n9136;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9138 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9139 = trap_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9140 = n9138 & n9139;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9141 = n9137 | n9140;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9142 = trap_ctrl[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9143 = csr[127]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9144 = n9142 & n9143;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9145 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9146 = trap_ctrl[43]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9147 = n9145 & n9146;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9148 = n9144 | n9147;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9149 = trap_ctrl[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9150 = csr[128]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9151 = n9149 & n9150;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9152 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9153 = trap_ctrl[44]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9154 = n9152 & n9153;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9155 = n9151 | n9154;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9156 = trap_ctrl[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9157 = csr[129]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9158 = n9156 & n9157;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9159 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9160 = trap_ctrl[45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9161 = n9159 & n9160;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9162 = n9158 | n9161;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9163 = trap_ctrl[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9164 = csr[130]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9165 = n9163 & n9164;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9166 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9167 = trap_ctrl[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9168 = n9166 & n9167;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9169 = n9165 | n9168;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9170 = trap_ctrl[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9171 = csr[131]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9172 = n9170 & n9171;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9173 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9174 = trap_ctrl[47]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9175 = n9173 & n9174;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9176 = n9172 | n9175;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9177 = trap_ctrl[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9178 = csr[132]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9179 = n9177 & n9178;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9180 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9181 = trap_ctrl[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9182 = n9180 & n9181;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9183 = n9179 | n9182;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9184 = trap_ctrl[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9185 = csr[133]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9186 = n9184 & n9185;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9187 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9188 = trap_ctrl[49]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9189 = n9187 & n9188;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9190 = n9186 | n9189;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9191 = trap_ctrl[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9192 = csr[134]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9193 = n9191 & n9192;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9194 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9195 = trap_ctrl[50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9196 = n9194 & n9195;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9197 = n9193 | n9196;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:64  */
  assign n9198 = trap_ctrl[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:97  */
  assign n9199 = csr[135]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:81  */
  assign n9200 = n9198 & n9199;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:116  */
  assign n9201 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:149  */
  assign n9202 = trap_ctrl[51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:128  */
  assign n9203 = n9201 & n9202;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1181:102  */
  assign n9204 = n9200 | n9203;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1185:54  */
  assign n9205 = debug_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1185:78  */
  assign n9206 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1185:111  */
  assign n9207 = trap_ctrl[52]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1185:90  */
  assign n9208 = n9206 & n9207;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1185:64  */
  assign n9209 = n9205 | n9208;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1186:54  */
  assign n9210 = debug_ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1186:78  */
  assign n9211 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1186:111  */
  assign n9212 = trap_ctrl[53]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1186:90  */
  assign n9213 = n9211 & n9212;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1186:64  */
  assign n9214 = n9210 | n9213;
  assign n9215 = {n9214, n9209, n9204, n9197, n9190, n9183, n9176, n9169, n9162, n9155, n9148, n9141, n9134, n9127, n9120, n9113, n9106, n9099, n9085, n9092, n9078, 1'b0, 1'b0, irq_fast_i, n9068, n9069, n9067};
  assign n9218 = {21'b000000000000000000000, 21'b000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1195:16  */
  assign n9222 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1200:31  */
  assign n9226 = trap_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1201:31  */
  assign n9228 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1202:31  */
  assign n9230 = trap_ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1203:31  */
  assign n9232 = trap_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1203:120  */
  assign n9234 = csr[136]; // extract
  assign n9240 = {n9234, n9234};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1203:102  */
  assign n9243 = {5'b00010, n9240};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1204:31  */
  assign n9244 = trap_ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1205:31  */
  assign n9246 = trap_ctrl[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1206:31  */
  assign n9248 = trap_ctrl[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1207:31  */
  assign n9250 = trap_ctrl[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1208:31  */
  assign n9252 = trap_ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1210:31  */
  assign n9254 = trap_ctrl[52]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1211:31  */
  assign n9256 = trap_ctrl[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1212:31  */
  assign n9258 = trap_ctrl[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1213:31  */
  assign n9260 = trap_ctrl[53]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1215:31  */
  assign n9262 = trap_ctrl[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1216:31  */
  assign n9264 = trap_ctrl[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1217:31  */
  assign n9266 = trap_ctrl[38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1218:31  */
  assign n9268 = trap_ctrl[39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1219:31  */
  assign n9270 = trap_ctrl[40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1220:31  */
  assign n9272 = trap_ctrl[41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1221:31  */
  assign n9274 = trap_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1222:31  */
  assign n9276 = trap_ctrl[43]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1223:31  */
  assign n9278 = trap_ctrl[44]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1224:31  */
  assign n9280 = trap_ctrl[45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1225:31  */
  assign n9282 = trap_ctrl[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1226:31  */
  assign n9284 = trap_ctrl[47]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1227:31  */
  assign n9286 = trap_ctrl[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1228:31  */
  assign n9288 = trap_ctrl[49]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1229:31  */
  assign n9290 = trap_ctrl[50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1230:31  */
  assign n9292 = trap_ctrl[51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1232:31  */
  assign n9294 = trap_ctrl[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1233:31  */
  assign n9296 = trap_ctrl[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1234:31  */
  assign n9298 = trap_ctrl[34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1234:7  */
  assign n9300 = n9298 ? 7'b1000111 : 7'b0000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1233:7  */
  assign n9301 = n9296 ? 7'b1000011 : n9300;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1232:7  */
  assign n9302 = n9294 ? 7'b1001011 : n9301;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1230:7  */
  assign n9303 = n9292 ? 7'b1011111 : n9302;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1229:7  */
  assign n9304 = n9290 ? 7'b1011110 : n9303;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1228:7  */
  assign n9305 = n9288 ? 7'b1011101 : n9304;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1227:7  */
  assign n9306 = n9286 ? 7'b1011100 : n9305;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1226:7  */
  assign n9307 = n9284 ? 7'b1011011 : n9306;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1225:7  */
  assign n9308 = n9282 ? 7'b1011010 : n9307;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1224:7  */
  assign n9309 = n9280 ? 7'b1011001 : n9308;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1223:7  */
  assign n9310 = n9278 ? 7'b1011000 : n9309;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1222:7  */
  assign n9311 = n9276 ? 7'b1010111 : n9310;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1221:7  */
  assign n9312 = n9274 ? 7'b1010110 : n9311;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1220:7  */
  assign n9313 = n9272 ? 7'b1010101 : n9312;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1219:7  */
  assign n9314 = n9270 ? 7'b1010100 : n9313;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1218:7  */
  assign n9315 = n9268 ? 7'b1010011 : n9314;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1217:7  */
  assign n9316 = n9266 ? 7'b1010010 : n9315;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1216:7  */
  assign n9317 = n9264 ? 7'b1010001 : n9316;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1215:7  */
  assign n9318 = n9262 ? 7'b1010000 : n9317;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1213:7  */
  assign n9319 = n9260 ? 7'b1100100 : n9318;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1212:7  */
  assign n9320 = n9258 ? 7'b0100001 : n9319;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1211:7  */
  assign n9321 = n9256 ? 7'b0100010 : n9320;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1210:7  */
  assign n9322 = n9254 ? 7'b1100011 : n9321;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1208:7  */
  assign n9323 = n9252 ? 7'b0000101 : n9322;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1207:7  */
  assign n9324 = n9250 ? 7'b0000111 : n9323;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1206:7  */
  assign n9325 = n9248 ? 7'b0000100 : n9324;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1205:7  */
  assign n9326 = n9246 ? 7'b0000110 : n9325;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1204:7  */
  assign n9327 = n9244 ? 7'b0000011 : n9326;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1203:7  */
  assign n9328 = n9232 ? n9243 : n9327;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1202:7  */
  assign n9329 = n9230 ? 7'b0000000 : n9328;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1201:7  */
  assign n9330 = n9228 ? 7'b0000010 : n9329;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1200:7  */
  assign n9331 = n9226 ? 7'b0000001 : n9330;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1240:31  */
  assign n9336 = exe_engine[100:69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1240:56  */
  assign n9337 = trap_ctrl[63]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1240:35  */
  assign n9338 = n9337 ? n9336 : n9339;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1240:102  */
  assign n9339 = exe_engine[68:37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1247:16  */
  assign n9341 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1252:21  */
  assign n9345 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1252:33  */
  assign n9346 = ~n9345;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1253:23  */
  assign n9347 = trap_ctrl[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9355 = trap_ctrl[56]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9357 = 1'b0 | n9355;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9359 = trap_ctrl[55]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9360 = n9357 | n9359;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9361 = trap_ctrl[54]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9362 = n9360 | n9361;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1253:39  */
  assign n9363 = n9347 | n9362;
  assign n9365 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1253:9  */
  assign n9366 = n9363 ? 1'b1 : n9365;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1257:23  */
  assign n9367 = trap_ctrl[97]; // extract
  assign n9369 = trap_ctrl[96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1257:9  */
  assign n9370 = n9367 ? 1'b0 : n9369;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1252:7  */
  assign n9371 = n9346 ? n9366 : n9370;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1262:22  */
  assign n9372 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1262:28  */
  assign n9374 = n9372 == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1264:24  */
  assign n9376 = trap_ctrl[97]; // extract
  assign n9378 = trap_ctrl[98]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1264:7  */
  assign n9379 = n9376 ? 1'b1 : n9378;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1262:7  */
  assign n9380 = n9374 ? 1'b0 : n9379;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9396 = trap_ctrl[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9398 = 1'b0 | n9396;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9400 = trap_ctrl[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9401 = n9398 | n9400;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9402 = trap_ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9403 = n9401 | n9402;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9404 = trap_ctrl[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9405 = n9403 | n9404;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9406 = trap_ctrl[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9407 = n9405 | n9406;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9408 = trap_ctrl[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9409 = n9407 | n9408;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9410 = trap_ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9411 = n9409 | n9410;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9412 = trap_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9413 = n9411 | n9412;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9414 = trap_ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9415 = n9413 | n9414;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9416 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9417 = n9415 | n9416;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9418 = trap_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9419 = n9417 | n9418;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1271:29  */
  assign n9420 = n9419 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1275:17  */
  assign n9423 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1275:23  */
  assign n9425 = n9423 == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9433 = trap_ctrl[51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9435 = 1'b0 | n9433;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9437 = trap_ctrl[50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9438 = n9435 | n9437;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9439 = trap_ctrl[49]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9440 = n9438 | n9439;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9441 = trap_ctrl[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9442 = n9440 | n9441;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9443 = trap_ctrl[47]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9444 = n9442 | n9443;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9445 = trap_ctrl[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9446 = n9444 | n9445;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9447 = trap_ctrl[45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9448 = n9446 | n9447;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9449 = trap_ctrl[44]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9450 = n9448 | n9449;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9451 = trap_ctrl[43]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9452 = n9450 | n9451;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9453 = trap_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9454 = n9452 | n9453;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9455 = trap_ctrl[41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9456 = n9454 | n9455;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9457 = trap_ctrl[40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9458 = n9456 | n9457;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9459 = trap_ctrl[39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9460 = n9458 | n9459;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9461 = trap_ctrl[38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9462 = n9460 | n9461;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9463 = trap_ctrl[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9464 = n9462 | n9463;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9465 = trap_ctrl[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9466 = n9464 | n9465;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9467 = trap_ctrl[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9468 = n9466 | n9467;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9469 = trap_ctrl[34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9470 = n9468 | n9469;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9471 = trap_ctrl[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9472 = n9470 | n9471;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1275:37  */
  assign n9473 = n9472 & n9425;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1277:11  */
  assign n9474 = csr[112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1277:38  */
  assign n9475 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1277:48  */
  assign n9476 = ~n9475;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1277:30  */
  assign n9477 = n9474 | n9476;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1276:80  */
  assign n9478 = n9477 & n9473;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1278:17  */
  assign n9479 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1278:21  */
  assign n9480 = ~n9479;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1277:66  */
  assign n9481 = n9480 & n9478;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1278:37  */
  assign n9482 = csr[324]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1278:47  */
  assign n9483 = ~n9482;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1278:28  */
  assign n9484 = n9483 & n9481;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1274:32  */
  assign n9485 = n9484 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1282:18  */
  assign n9488 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1282:24  */
  assign n9490 = n9488 == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1282:53  */
  assign n9491 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1282:59  */
  assign n9493 = n9491 == 4'b1000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1282:38  */
  assign n9494 = n9490 | n9493;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1283:23  */
  assign n9495 = trap_ctrl[52]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1282:75  */
  assign n9496 = n9495 & n9494;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1281:32  */
  assign n9497 = n9496 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1287:18  */
  assign n9500 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1287:24  */
  assign n9502 = n9500 == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1288:18  */
  assign n9503 = trap_ctrl[98]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1288:53  */
  assign n9504 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1288:59  */
  assign n9506 = n9504 == 4'b1000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1288:37  */
  assign n9507 = n9506 & n9503;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1287:38  */
  assign n9508 = n9502 | n9507;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1289:23  */
  assign n9509 = trap_ctrl[53]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1288:76  */
  assign n9510 = n9509 & n9508;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1286:32  */
  assign n9511 = n9510 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1296:16  */
  assign n9514 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1299:22  */
  assign n9516 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1299:28  */
  assign n9518 = n9516 == 4'b0100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1300:15  */
  assign n9519 = ipb[73:72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1300:20  */
  assign n9521 = n9519 != 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1299:40  */
  assign n9522 = n9521 & n9518;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1301:21  */
  assign n9523 = trap_ctrl[100]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1301:28  */
  assign n9524 = ~n9523;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1300:29  */
  assign n9525 = n9524 & n9522;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1299:7  */
  assign n9528 = n9525 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9540 = trap_ctrl[53]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9542 = 1'b0 | n9540;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9544 = trap_ctrl[52]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9545 = n9542 | n9544;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9546 = trap_ctrl[51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9547 = n9545 | n9546;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9548 = trap_ctrl[50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9549 = n9547 | n9548;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9550 = trap_ctrl[49]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9551 = n9549 | n9550;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9552 = trap_ctrl[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9553 = n9551 | n9552;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9554 = trap_ctrl[47]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9555 = n9553 | n9554;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9556 = trap_ctrl[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9557 = n9555 | n9556;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9558 = trap_ctrl[45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9559 = n9557 | n9558;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9560 = trap_ctrl[44]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9561 = n9559 | n9560;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9562 = trap_ctrl[43]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9563 = n9561 | n9562;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9564 = trap_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9565 = n9563 | n9564;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9566 = trap_ctrl[41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9567 = n9565 | n9566;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9568 = trap_ctrl[40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9569 = n9567 | n9568;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9570 = trap_ctrl[39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9571 = n9569 | n9570;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9572 = trap_ctrl[38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9573 = n9571 | n9572;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9574 = trap_ctrl[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9575 = n9573 | n9574;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9576 = trap_ctrl[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9577 = n9575 | n9576;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9578 = trap_ctrl[35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9579 = n9577 | n9578;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9580 = trap_ctrl[34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9581 = n9579 | n9580;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n9582 = trap_ctrl[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n9583 = n9581 | n9582;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1310:68  */
  assign n9584 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1310:54  */
  assign n9585 = n9583 | n9584;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1310:79  */
  assign n9586 = csr[324]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1310:72  */
  assign n9587 = n9585 | n9586;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1321:16  */
  assign n9589 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1324:18  */
  assign n9593 = opcode == 7'b1110011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1325:34  */
  assign n9594 = exe_engine[35:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1333:46  */
  assign n9601 = exe_engine[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1333:67  */
  assign n9602 = ~n9601;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1333:27  */
  assign n9603 = n9602 ? rf_rs1_i : n9606;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1333:113  */
  assign n9604 = exe_engine[23:19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1333:98  */
  assign n9606 = {27'b000000000000000000000000000, n9604};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1336:21  */
  assign n9607 = exe_engine[17:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1337:9  */
  assign n9608 = csr[111:80]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1337:28  */
  assign n9609 = csr[47:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1337:15  */
  assign n9610 = n9608 | n9609;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1337:37  */
  assign n9612 = n9607 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1338:9  */
  assign n9613 = csr[111:80]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1338:28  */
  assign n9614 = csr[47:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1338:20  */
  assign n9615 = ~n9614;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1338:15  */
  assign n9616 = n9613 & n9615;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1338:37  */
  assign n9618 = n9607 == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1339:9  */
  assign n9619 = csr[47:16]; // extract
  assign n9620 = {n9618, n9612};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1336:3  */
  always @*
    case (n9620)
      2'b10: n9621 = n9616;
      2'b01: n9621 = n9610;
      default: n9621 = n9619;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1344:23  */
  assign n9622 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1345:23  */
  assign n9623 = csr[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1346:23  */
  assign n9624 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1347:23  */
  assign n9625 = csr[79:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1354:16  */
  assign n9627 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1389:21  */
  assign n9660 = csr[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1389:54  */
  assign n9661 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1389:33  */
  assign n9662 = ~n9661;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1389:28  */
  assign n9663 = n9660 & n9662;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:15  */
  assign n9664 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1401:17  */
  assign n9665 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1401:22  */
  assign n9667 = n9665 == 12'b001100000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1402:40  */
  assign n9668 = csr[51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1403:40  */
  assign n9669 = csr[55]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1405:42  */
  assign n9670 = csr[59]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1405:59  */
  assign n9671 = csr[60]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1405:47  */
  assign n9672 = n9670 | n9671;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1406:42  */
  assign n9673 = csr[65]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1407:42  */
  assign n9674 = csr[69]; // extract
  assign n9675 = {n9674, n9673, n9672, n9669, n9668};
  assign n9676 = csr[116:112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1401:9  */
  assign n9677 = n9667 ? n9675 : n9676;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1412:17  */
  assign n9678 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1412:22  */
  assign n9680 = n9678 == 12'b001100000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1413:36  */
  assign n9681 = csr[51]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1414:36  */
  assign n9682 = csr[55]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1415:36  */
  assign n9683 = csr[59]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1416:36  */
  assign n9684 = csr[79:64]; // extract
  assign n9685 = {n9684, n9682, n9683, n9681};
  assign n9686 = csr[135:117]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1412:9  */
  assign n9687 = n9680 ? n9685 : n9686;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1420:17  */
  assign n9688 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1420:22  */
  assign n9690 = n9688 == 12'b001100000101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1421:33  */
  assign n9691 = csr[79:50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1421:51  */
  assign n9693 = {n9691, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1421:68  */
  assign n9694 = csr[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1421:57  */
  assign n9695 = {n9693, n9694};
  assign n9696 = csr[207:176]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1420:9  */
  assign n9697 = n9690 ? n9695 : n9696;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1425:17  */
  assign n9698 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1425:22  */
  assign n9700 = n9698 == 12'b001100000110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1425:42  */
  assign n9702 = 1'b1 & n9700;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1425:58  */
  assign n9704 = 1'b1 & n9702;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1426:41  */
  assign n9705 = csr[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1427:41  */
  assign n9706 = csr[50]; // extract
  assign n9707 = {n9706, n9705};
  assign n9708 = csr[305:304]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1425:9  */
  assign n9709 = n9704 ? n9707 : n9708;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1435:17  */
  assign n9710 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1435:22  */
  assign n9712 = n9710 == 12'b001101000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1436:31  */
  assign n9713 = csr[79:48]; // extract
  assign n9714 = csr[303:272]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1435:9  */
  assign n9715 = n9712 ? n9713 : n9714;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1440:17  */
  assign n9716 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1440:22  */
  assign n9718 = n9716 == 12'b001101000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1441:32  */
  assign n9719 = csr[79:49]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1441:50  */
  assign n9721 = {n9719, 1'b0};
  assign n9722 = csr[169:138]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1440:9  */
  assign n9723 = n9718 ? n9721 : n9722;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1448:17  */
  assign n9724 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1448:22  */
  assign n9726 = n9724 == 12'b001101000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1449:34  */
  assign n9727 = csr[79]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1449:50  */
  assign n9728 = csr[52:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1449:39  */
  assign n9729 = {n9727, n9728};
  assign n9730 = csr[175:170]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1448:9  */
  assign n9731 = n9726 ? n9729 : n9730;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1457:17  */
  assign n9732 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1457:22  */
  assign n9734 = n9732 == 12'b001100100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1459:46  */
  assign n9735 = csr[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1460:46  */
  assign n9736 = csr[50]; // extract
  assign n9737 = csr[306]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1457:9  */
  assign n9738 = n9734 ? n9735 : n9737;
  assign n9739 = csr[308]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9740 = n9944 ? n9736 : n9739;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1472:17  */
  assign n9741 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1472:22  */
  assign n9743 = n9741 == 12'b011110110000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1472:36  */
  assign n9745 = 1'b1 & n9743;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1473:40  */
  assign n9746 = csr[63]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1474:40  */
  assign n9747 = csr[50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1476:42  */
  assign n9748 = csr[60]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1477:42  */
  assign n9749 = csr[49]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1477:58  */
  assign n9750 = csr[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1477:46  */
  assign n9751 = n9749 | n9750;
  assign n9752 = {n9751, n9747, n9748, n9746};
  assign n9753 = csr[325:322]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1472:9  */
  assign n9754 = n9745 ? n9752 : n9753;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1482:17  */
  assign n9755 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1482:22  */
  assign n9757 = n9755 == 12'b011110110001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1482:35  */
  assign n9759 = 1'b1 & n9757;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1483:31  */
  assign n9760 = csr[79:49]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1483:49  */
  assign n9762 = {n9760, 1'b0};
  assign n9763 = csr[392:361]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1482:9  */
  assign n9764 = n9759 ? n9762 : n9763;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1490:17  */
  assign n9765 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1490:22  */
  assign n9767 = n9765 == 12'b011110110010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1490:41  */
  assign n9769 = 1'b1 & n9767;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1491:32  */
  assign n9770 = csr[79:48]; // extract
  assign n9771 = csr[424:393]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1490:9  */
  assign n9772 = n9769 ? n9770 : n9771;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1499:17  */
  assign n9773 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1499:22  */
  assign n9775 = n9773 == 12'b011110100001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1499:38  */
  assign n9777 = 1'b1 & n9775;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1500:19  */
  assign n9778 = csr[427]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1500:32  */
  assign n9779 = ~n9778;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1500:54  */
  assign n9780 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1500:39  */
  assign n9781 = n9779 | n9780;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1501:44  */
  assign n9782 = csr[50]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1502:44  */
  assign n9783 = csr[60]; // extract
  assign n9784 = {n9783, n9782};
  assign n9785 = csr[426:425]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1500:11  */
  assign n9786 = n9781 ? n9784 : n9785;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1504:26  */
  assign n9787 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1505:42  */
  assign n9788 = csr[75]; // extract
  assign n9789 = csr[427]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1504:11  */
  assign n9790 = n9787 ? n9788 : n9789;
  assign n9791 = {n9790, n9786};
  assign n9792 = csr[427:425]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1499:9  */
  assign n9793 = n9777 ? n9791 : n9792;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1510:17  */
  assign n9794 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1510:22  */
  assign n9796 = n9794 == 12'b011110100010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1510:38  */
  assign n9798 = 1'b1 & n9796;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1511:19  */
  assign n9799 = csr[427]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1511:32  */
  assign n9800 = ~n9799;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1511:54  */
  assign n9801 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1511:39  */
  assign n9802 = n9800 | n9801;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1512:36  */
  assign n9803 = csr[79:49]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1512:54  */
  assign n9805 = {n9803, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1510:9  */
  assign n9809 = n9802 & n9798;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:24  */
  assign n9810 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1522:54  */
  assign n9811 = trap_ctrl[62]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1522:58  */
  assign n9812 = ~n9811;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1522:81  */
  assign n9813 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1522:85  */
  assign n9814 = ~n9813;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1522:65  */
  assign n9815 = n9814 & n9812;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1522:34  */
  assign n9817 = 1'b0 | n9815;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1523:40  */
  assign n9818 = trap_ctrl[63]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1523:80  */
  assign n9819 = trap_ctrl[61:57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1523:63  */
  assign n9820 = {n9818, n9819};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1524:38  */
  assign n9821 = trap_ctrl[95:65]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1524:56  */
  assign n9823 = {n9821, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1526:30  */
  assign n9824 = trap_ctrl[63]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1526:34  */
  assign n9825 = ~n9824;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1526:61  */
  assign n9826 = trap_ctrl[59]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1526:41  */
  assign n9827 = n9826 & n9825;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1526:11  */
  assign n9829 = n9827 ? lsu_mar_i : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1532:30  */
  assign n9830 = trap_ctrl[63]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1532:34  */
  assign n9831 = ~n9830;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1534:28  */
  assign n9833 = exe_engine[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1534:38  */
  assign n9835 = 1'b1 & n9833;
  assign n9837 = exe_engine[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1534:13  */
  assign n9838 = n9835 ? 1'b0 : n9837;
  assign n9839 = exe_engine[35:6]; // extract
  assign n9840 = exe_engine[4]; // extract
  assign n9842 = {n9839, n9838, n9840};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1532:11  */
  assign n9843 = n9831 ? n9842 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1543:35  */
  assign n9846 = csr[112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1544:35  */
  assign n9847 = csr[136]; // extract
  assign n9848 = {n9847, n9846, 1'b0};
  assign n9849 = {n9820, n9823};
  assign n9850 = {n9843, n9829};
  assign n9851 = csr[114:112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1522:9  */
  assign n9852 = n9817 ? n9848 : n9851;
  assign n9853 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1522:9  */
  assign n9854 = n9817 ? 1'b1 : n9853;
  assign n9855 = csr[175:138]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9856 = n9915 ? n9849 : n9855;
  assign n9857 = csr[271:208]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9858 = n9917 ? n9850 : n9857;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1548:48  */
  assign n9859 = trap_ctrl[62]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1548:28  */
  assign n9861 = n9859 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1548:75  */
  assign n9862 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1548:79  */
  assign n9863 = ~n9862;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1548:59  */
  assign n9864 = n9863 & n9861;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1549:44  */
  assign n9865 = trap_ctrl[59:57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1550:33  */
  assign n9866 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1551:42  */
  assign n9867 = trap_ctrl[95:65]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1551:60  */
  assign n9869 = {n9867, 1'b0};
  assign n9870 = {n9865, n9866};
  assign n9871 = csr[328:325]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9872 = n9919 ? n9870 : n9871;
  assign n9873 = csr[392:361]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9874 = n9921 ? n9869 : n9873;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1557:24  */
  assign n9875 = trap_ctrl[99]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1560:44  */
  assign n9876 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1560:28  */
  assign n9878 = n9876 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1562:34  */
  assign n9879 = csr[325]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1563:21  */
  assign n9880 = csr[325]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1563:30  */
  assign n9882 = n9880 != 1'b1;
  assign n9884 = csr[115]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1563:13  */
  assign n9885 = n9882 ? 1'b0 : n9884;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1570:36  */
  assign n9886 = csr[114]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1572:21  */
  assign n9888 = csr[114]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1572:33  */
  assign n9890 = n9888 != 1'b1;
  assign n9892 = csr[115]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1572:13  */
  assign n9893 = n9890 ? 1'b0 : n9892;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1576:35  */
  assign n9894 = csr[113]; // extract
  assign n9896 = {n9893, 1'b0, 1'b1, n9894};
  assign n9897 = n9896[2:0]; // extract
  assign n9898 = csr[114:112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1560:9  */
  assign n9899 = n9878 ? n9898 : n9897;
  assign n9900 = n9896[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1560:9  */
  assign n9901 = n9878 ? n9885 : n9900;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1560:9  */
  assign n9902 = n9878 ? n9879 : n9886;
  assign n9903 = {n9901, n9899};
  assign n9904 = csr[115:112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1557:7  */
  assign n9905 = n9875 ? n9903 : n9904;
  assign n9906 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1557:7  */
  assign n9907 = n9875 ? n9902 : n9906;
  assign n9908 = n9905[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9909 = n9810 ? n9852 : n9908;
  assign n9910 = n9905[3]; // extract
  assign n9911 = csr[115]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9912 = n9810 ? n9911 : n9910;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9913 = n9810 ? n9854 : n9907;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9915 = n9817 & n9810;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9917 = n9817 & n9810;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9919 = n9864 & n9810;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1519:7  */
  assign n9921 = n9864 & n9810;
  assign n9922 = {n9912, n9909};
  assign n9923 = {n9687, n9677};
  assign n9924 = {n9697, n9731, n9723};
  assign n9925 = {n9738, n9709, n9715};
  assign n9926 = {n9793, n9772, n9764};
  assign n9927 = n9923[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9928 = n9664 ? n9927 : n9922;
  assign n9929 = n9923[23:4]; // extract
  assign n9930 = csr[135:116]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9931 = n9664 ? n9929 : n9930;
  assign n9932 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9933 = n9664 ? n9932 : n9913;
  assign n9934 = n9924[37:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9935 = n9664 ? n9934 : n9856;
  assign n9936 = n9924[69:38]; // extract
  assign n9937 = csr[207:176]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9938 = n9664 ? n9936 : n9937;
  assign n9939 = csr[271:208]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9940 = n9664 ? n9939 : n9858;
  assign n9941 = csr[306:272]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9942 = n9664 ? n9925 : n9941;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9944 = n9734 & n9664;
  assign n9945 = n9754[2:0]; // extract
  assign n9946 = csr[324:322]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9947 = n9664 ? n9945 : n9946;
  assign n9948 = n9872[0]; // extract
  assign n9949 = n9754[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9950 = n9664 ? n9949 : n9948;
  assign n9951 = n9872[3:1]; // extract
  assign n9952 = csr[328:326]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9953 = n9664 ? n9952 : n9951;
  assign n9954 = n9926[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9955 = n9664 ? n9954 : n9874;
  assign n9956 = n9926[66:32]; // extract
  assign n9957 = csr[427:393]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9958 = n9664 ? n9956 : n9957;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1394:7  */
  assign n9960 = n9809 & n9664;
  assign n9963 = {n9933, n9931, n9928};
  assign n9964 = {n9953, n9950, n9947, 13'b0000000000000, n9740, 1'b0, n9942, n9940, n9938, n9935};
  assign n9965 = {n9958, n9955};
  assign n9976 = {1'b1, 16'b0000000000000000, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0};
  assign n9977 = {3'b000, 1'b0, 1'b0, 1'b0, 1'b0, 16'b0000000000000000, 1'b0, 1'b0, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 6'b000000, 32'b00000000000000000000000000000000};
  assign n9978 = {1'b0, 1'b0, 1'b0, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1640:55  */
  assign n9986 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1640:38  */
  assign n9987 = n9986 ? 1'b1 : n9988;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1640:75  */
  assign n9988 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1647:16  */
  assign n9990 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1651:24  */
  assign n9994 = csr[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1651:57  */
  assign n9995 = trap_ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1651:36  */
  assign n9996 = ~n9995;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1651:31  */
  assign n9997 = n9994 & n9996;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1653:15  */
  assign n9999 = csr[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:18  */
  assign n10000 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1659:11  */
  assign n10002 = n10000 == 12'b000000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1659:29  */
  assign n10004 = n10000 == 12'b000000000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1659:29  */
  assign n10005 = n10002 | n10004;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1659:41  */
  assign n10007 = n10000 == 12'b000000000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1659:41  */
  assign n10008 = n10005 | n10007;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1667:11  */
  assign n10010 = n10000 == 12'b100000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1667:30  */
  assign n10012 = n10000 == 12'b100000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1667:30  */
  assign n10013 = n10010 | n10012;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1667:46  */
  assign n10015 = n10000 == 12'b100000000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1667:46  */
  assign n10016 = n10013 | n10015;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1667:62  */
  assign n10018 = n10000 == 12'b100000000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1667:62  */
  assign n10019 = n10016 | n10018;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1675:11  */
  assign n10021 = n10000 == 12'b101111000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1675:32  */
  assign n10023 = n10000 == 12'b101111000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1675:32  */
  assign n10024 = n10021 | n10023;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1682:34  */
  assign n10025 = csr[112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1683:34  */
  assign n10026 = csr[113]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1684:55  */
  assign n10027 = csr[114]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1684:55  */
  assign n10028 = csr[114]; // extract
  assign n10029 = {n10027, n10028};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1685:34  */
  assign n10030 = csr[115]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1686:34  */
  assign n10031 = csr[116]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1686:45  */
  assign n10034 = n10031 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1681:11  */
  assign n10036 = n10000 == 12'b001100000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1690:11  */
  assign n10052 = n10000 == 12'b001100000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1701:34  */
  assign n10053 = csr[117]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1702:34  */
  assign n10054 = csr[119]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1703:34  */
  assign n10055 = csr[118]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1704:44  */
  assign n10056 = csr[135:120]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1700:11  */
  assign n10058 = n10000 == 12'b001100000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1707:30  */
  assign n10059 = csr[207:176]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1706:11  */
  assign n10061 = n10000 == 12'b001100000101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1711:35  */
  assign n10062 = csr[304]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1712:35  */
  assign n10063 = csr[305]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1709:11  */
  assign n10065 = n10000 == 12'b001100000110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1725:30  */
  assign n10066 = csr[303:272]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1724:11  */
  assign n10068 = n10000 == 12'b001101000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1728:34  */
  assign n10069 = csr[169:139]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1728:52  */
  assign n10071 = {n10069, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1727:11  */
  assign n10073 = n10000 == 12'b001101000001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1731:48  */
  assign n10074 = csr[175]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1732:48  */
  assign n10075 = csr[174:170]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1730:11  */
  assign n10077 = n10000 == 12'b001101000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1735:30  */
  assign n10078 = csr[239:208]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1734:11  */
  assign n10080 = n10000 == 12'b001101000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1738:57  */
  assign n10081 = trap_ctrl[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1739:57  */
  assign n10082 = trap_ctrl[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1740:57  */
  assign n10083 = trap_ctrl[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1741:57  */
  assign n10084 = trap_ctrl[30:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1737:11  */
  assign n10086 = n10000 == 12'b001101000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1744:30  */
  assign n10087 = csr[271:240]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1743:11  */
  assign n10089 = n10000 == 12'b001101001010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:11  */
  assign n10091 = n10000 == 12'b001110100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:32  */
  assign n10093 = n10000 == 12'b001110100001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:32  */
  assign n10094 = n10091 | n10093;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:50  */
  assign n10096 = n10000 == 12'b001110100010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:50  */
  assign n10097 = n10094 | n10096;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:68  */
  assign n10099 = n10000 == 12'b001110100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:68  */
  assign n10100 = n10097 | n10099;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:86  */
  assign n10102 = n10000 == 12'b001110110000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1749:86  */
  assign n10103 = n10100 | n10102;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1750:32  */
  assign n10105 = n10000 == 12'b001110110001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1750:32  */
  assign n10106 = n10103 | n10105;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1750:50  */
  assign n10108 = n10000 == 12'b001110110010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1750:50  */
  assign n10109 = n10106 | n10108;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1750:68  */
  assign n10111 = n10000 == 12'b001110110011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1750:68  */
  assign n10112 = n10109 | n10111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1750:86  */
  assign n10114 = n10000 == 12'b001110110100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1750:86  */
  assign n10115 = n10112 | n10114;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1751:32  */
  assign n10117 = n10000 == 12'b001110110101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1751:32  */
  assign n10118 = n10115 | n10117;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1751:50  */
  assign n10120 = n10000 == 12'b001110110110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1751:50  */
  assign n10121 = n10118 | n10120;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1751:68  */
  assign n10123 = n10000 == 12'b001110110111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1751:68  */
  assign n10124 = n10121 | n10123;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1751:86  */
  assign n10126 = n10000 == 12'b001110111000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1751:86  */
  assign n10127 = n10124 | n10126;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1752:32  */
  assign n10129 = n10000 == 12'b001110111001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1752:32  */
  assign n10130 = n10127 | n10129;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1752:50  */
  assign n10132 = n10000 == 12'b001110111010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1752:50  */
  assign n10133 = n10130 | n10132;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1752:68  */
  assign n10135 = n10000 == 12'b001110111011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1752:68  */
  assign n10136 = n10133 | n10135;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1752:86  */
  assign n10138 = n10000 == 12'b001110111100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1752:86  */
  assign n10139 = n10136 | n10138;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1753:32  */
  assign n10141 = n10000 == 12'b001110111101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1753:32  */
  assign n10142 = n10139 | n10141;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1753:50  */
  assign n10144 = n10000 == 12'b001110111110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1753:50  */
  assign n10145 = n10142 | n10144;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1753:68  */
  assign n10147 = n10000 == 12'b001110111111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1753:68  */
  assign n10148 = n10145 | n10147;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1763:48  */
  assign n10149 = csr[306]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1764:48  */
  assign n10150 = csr[308]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1761:11  */
  assign n10152 = n10000 == 12'b001100100000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1773:11  */
  assign n10154 = n10000 == 12'b001100100011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1774:11  */
  assign n10156 = n10000 == 12'b001100100100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1775:11  */
  assign n10158 = n10000 == 12'b001100100101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1776:11  */
  assign n10160 = n10000 == 12'b001100100110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1777:11  */
  assign n10162 = n10000 == 12'b001100100111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1778:11  */
  assign n10164 = n10000 == 12'b001100101000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1779:11  */
  assign n10166 = n10000 == 12'b001100101001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1780:11  */
  assign n10168 = n10000 == 12'b001100101010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1781:11  */
  assign n10170 = n10000 == 12'b001100101011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1782:11  */
  assign n10172 = n10000 == 12'b001100101100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1783:11  */
  assign n10174 = n10000 == 12'b001100101101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1784:11  */
  assign n10176 = n10000 == 12'b001100101110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1785:11  */
  assign n10178 = n10000 == 12'b001100101111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1791:97  */
  assign n10179 = cnt_lo_rd[95:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1791:11  */
  assign n10181 = n10000 == 12'b101100000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1791:31  */
  assign n10183 = n10000 == 12'b110000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1791:31  */
  assign n10184 = n10181 | n10183;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1792:97  */
  assign n10185 = cnt_lo_rd[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1792:11  */
  assign n10187 = n10000 == 12'b101100000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1792:31  */
  assign n10189 = n10000 == 12'b110000000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1792:31  */
  assign n10190 = n10187 | n10189;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1793:11  */
  assign n10192 = n10000 == 12'b101100000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1794:11  */
  assign n10194 = n10000 == 12'b101100000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1795:11  */
  assign n10196 = n10000 == 12'b101100000101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1796:11  */
  assign n10198 = n10000 == 12'b101100000110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1797:11  */
  assign n10200 = n10000 == 12'b101100000111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1798:11  */
  assign n10202 = n10000 == 12'b101100001000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1799:11  */
  assign n10204 = n10000 == 12'b101100001001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1800:11  */
  assign n10206 = n10000 == 12'b101100001010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1801:11  */
  assign n10208 = n10000 == 12'b101100001011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1802:11  */
  assign n10210 = n10000 == 12'b101100001100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1803:11  */
  assign n10212 = n10000 == 12'b101100001101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1804:11  */
  assign n10214 = n10000 == 12'b101100001110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1805:11  */
  assign n10216 = n10000 == 12'b101100001111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1808:99  */
  assign n10217 = cnt_hi_rd[95:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1808:11  */
  assign n10219 = n10000 == 12'b101110000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1808:32  */
  assign n10221 = n10000 == 12'b110010000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1808:32  */
  assign n10222 = n10219 | n10221;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1809:99  */
  assign n10223 = cnt_hi_rd[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1809:11  */
  assign n10225 = n10000 == 12'b101110000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1809:32  */
  assign n10227 = n10000 == 12'b110010000010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1809:32  */
  assign n10228 = n10225 | n10227;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1810:11  */
  assign n10230 = n10000 == 12'b101110000011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1811:11  */
  assign n10232 = n10000 == 12'b101110000100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1812:11  */
  assign n10234 = n10000 == 12'b101110000101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1813:11  */
  assign n10236 = n10000 == 12'b101110000110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1814:11  */
  assign n10238 = n10000 == 12'b101110000111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1815:11  */
  assign n10240 = n10000 == 12'b101110001000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1816:11  */
  assign n10242 = n10000 == 12'b101110001001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1817:11  */
  assign n10244 = n10000 == 12'b101110001010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1818:11  */
  assign n10246 = n10000 == 12'b101110001011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1819:11  */
  assign n10248 = n10000 == 12'b101110001100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1820:11  */
  assign n10250 = n10000 == 12'b101110001101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1821:11  */
  assign n10252 = n10000 == 12'b101110001110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1822:11  */
  assign n10254 = n10000 == 12'b101110001111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1827:11  */
  assign n10257 = n10000 == 12'b111100010001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1828:11  */
  assign n10260 = n10000 == 12'b111100010010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1829:11  */
  assign n10263 = n10000 == 12'b111100010011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1830:11  */
  assign n10266 = n10000 == 12'b111100010100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1836:76  */
  assign n10267 = csr[360:329]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1836:11  */
  assign n10269 = n10000 == 12'b011110110000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1837:76  */
  assign n10270 = csr[392:361]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1837:11  */
  assign n10272 = n10000 == 12'b011110110001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1838:76  */
  assign n10273 = csr[424:393]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1838:11  */
  assign n10275 = n10000 == 12'b011110110010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1844:75  */
  assign n10276 = csr[459:428]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1844:11  */
  assign n10278 = n10000 == 12'b011110100001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1845:75  */
  assign n10279 = csr[491:460]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1845:11  */
  assign n10281 = n10000 == 12'b011110100010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1846:11  */
  assign n10284 = n10000 == 12'b011110100100;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1852:11  */
  assign n10347 = n10000 == 12'b111111000000;
  assign n10348 = {n10347, n10284, n10281, n10278, n10275, n10272, n10269, n10266, n10263, n10260, n10257, n10254, n10252, n10250, n10248, n10246, n10244, n10242, n10240, n10238, n10236, n10234, n10232, n10230, n10228, n10222, n10216, n10214, n10212, n10210, n10208, n10206, n10204, n10202, n10200, n10198, n10196, n10194, n10192, n10190, n10184, n10178, n10176, n10174, n10172, n10170, n10168, n10166, n10164, n10162, n10160, n10158, n10156, n10154, n10152, n10148, n10089, n10086, n10080, n10077, n10073, n10068, n10065, n10061, n10058, n10052, n10036, n10024, n10019, n10008};
  assign n10349 = xcsr_rdata_i[0]; // extract
  assign n10350 = n10059[0]; // extract
  assign n10351 = n10066[0]; // extract
  assign n10352 = n10071[0]; // extract
  assign n10353 = n10075[0]; // extract
  assign n10354 = n10078[0]; // extract
  assign n10355 = n10087[0]; // extract
  assign n10356 = n10179[0]; // extract
  assign n10357 = n10185[0]; // extract
  assign n10358 = n10217[0]; // extract
  assign n10359 = n10223[0]; // extract
  assign n10360 = n10255[0]; // extract
  assign n10361 = n10258[0]; // extract
  assign n10362 = n10261[0]; // extract
  assign n10363 = n10264[0]; // extract
  assign n10364 = n10267[0]; // extract
  assign n10365 = n10270[0]; // extract
  assign n10366 = n10273[0]; // extract
  assign n10367 = n10276[0]; // extract
  assign n10368 = n10279[0]; // extract
  assign n10369 = n10282[0]; // extract
  assign n10370 = n9998[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10371 = 1'b1;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10371 = n10369;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10371 = n10368;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10371 = n10367;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10371 = n10366;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10371 = n10365;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10371 = n10364;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10371 = n10363;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10371 = n10362;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10371 = n10361;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10371 = n10360;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10371 = n10359;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10371 = n10358;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10371 = n10357;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10371 = n10356;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10371 = n10149;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10371 = n10355;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10371 = n10354;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10371 = n10353;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10371 = n10352;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10371 = n10351;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10371 = n10062;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10371 = n10350;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10371 = n10349;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10371 = n10370;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10371 = n10370;
      default: n10371 = n10370;
    endcase
  assign n10372 = xcsr_rdata_i[1]; // extract
  assign n10373 = n10059[1]; // extract
  assign n10374 = n10066[1]; // extract
  assign n10375 = n10071[1]; // extract
  assign n10376 = n10075[1]; // extract
  assign n10377 = n10078[1]; // extract
  assign n10378 = n10087[1]; // extract
  assign n10379 = n10179[1]; // extract
  assign n10380 = n10185[1]; // extract
  assign n10381 = n10217[1]; // extract
  assign n10382 = n10223[1]; // extract
  assign n10383 = n10255[1]; // extract
  assign n10384 = n10258[1]; // extract
  assign n10385 = n10261[1]; // extract
  assign n10386 = n10264[1]; // extract
  assign n10387 = n10267[1]; // extract
  assign n10388 = n10270[1]; // extract
  assign n10389 = n10273[1]; // extract
  assign n10390 = n10276[1]; // extract
  assign n10391 = n10279[1]; // extract
  assign n10392 = n10282[1]; // extract
  assign n10393 = n9998[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10394 = 1'b1;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10394 = n10392;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10394 = n10391;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10394 = n10390;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10394 = n10389;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10394 = n10388;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10394 = n10387;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10394 = n10386;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10394 = n10385;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10394 = n10384;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10394 = n10383;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10394 = n10382;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10394 = n10381;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10394 = n10380;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10394 = n10379;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10394 = n10378;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10394 = n10377;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10394 = n10376;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10394 = n10375;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10394 = n10374;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10394 = n10373;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10394 = 1'b0;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10394 = n10372;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10394 = n10393;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10394 = n10393;
      default: n10394 = n10393;
    endcase
  assign n10395 = xcsr_rdata_i[2]; // extract
  assign n10396 = n10059[2]; // extract
  assign n10397 = n10066[2]; // extract
  assign n10398 = n10071[2]; // extract
  assign n10399 = n10075[2]; // extract
  assign n10400 = n10078[2]; // extract
  assign n10401 = n10087[2]; // extract
  assign n10402 = n10179[2]; // extract
  assign n10403 = n10185[2]; // extract
  assign n10404 = n10217[2]; // extract
  assign n10405 = n10223[2]; // extract
  assign n10406 = n10255[2]; // extract
  assign n10407 = n10258[2]; // extract
  assign n10408 = n10261[2]; // extract
  assign n10409 = n10264[2]; // extract
  assign n10410 = n10267[2]; // extract
  assign n10411 = n10270[2]; // extract
  assign n10412 = n10273[2]; // extract
  assign n10413 = n10276[2]; // extract
  assign n10414 = n10279[2]; // extract
  assign n10415 = n10282[2]; // extract
  assign n10416 = n9998[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10417 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10417 = n10415;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10417 = n10414;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10417 = n10413;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10417 = n10412;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10417 = n10411;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10417 = n10410;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10417 = n10409;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10417 = n10408;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10417 = n10407;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10417 = n10406;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10417 = n10405;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10417 = n10404;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10417 = n10403;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10417 = n10402;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10417 = n10150;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10417 = n10401;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10417 = n10400;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10417 = n10399;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10417 = n10398;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10417 = n10397;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10417 = n10063;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10417 = n10396;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10417 = 1'b1;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10417 = n10395;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10417 = n10416;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10417 = n10416;
      default: n10417 = n10416;
    endcase
  assign n10418 = xcsr_rdata_i[3]; // extract
  assign n10419 = n10059[3]; // extract
  assign n10420 = n10066[3]; // extract
  assign n10421 = n10071[3]; // extract
  assign n10422 = n10075[3]; // extract
  assign n10423 = n10078[3]; // extract
  assign n10424 = n10087[3]; // extract
  assign n10425 = n10179[3]; // extract
  assign n10426 = n10185[3]; // extract
  assign n10427 = n10217[3]; // extract
  assign n10428 = n10223[3]; // extract
  assign n10429 = n10255[3]; // extract
  assign n10430 = n10258[3]; // extract
  assign n10431 = n10261[3]; // extract
  assign n10432 = n10264[3]; // extract
  assign n10433 = n10267[3]; // extract
  assign n10434 = n10270[3]; // extract
  assign n10435 = n10273[3]; // extract
  assign n10436 = n10276[3]; // extract
  assign n10437 = n10279[3]; // extract
  assign n10438 = n10282[3]; // extract
  assign n10439 = n9998[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10440 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10440 = n10438;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10440 = n10437;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10440 = n10436;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10440 = n10435;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10440 = n10434;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10440 = n10433;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10440 = n10432;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10440 = n10431;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10440 = n10430;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10440 = n10429;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10440 = n10428;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10440 = n10427;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10440 = n10426;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10440 = n10425;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10440 = n10424;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10440 = n10081;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10440 = n10423;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10440 = n10422;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10440 = n10421;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10440 = n10420;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10440 = n10419;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10440 = n10053;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10440 = n10025;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10440 = n10418;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10440 = n10439;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10440 = n10439;
      default: n10440 = n10439;
    endcase
  assign n10441 = xcsr_rdata_i[4]; // extract
  assign n10442 = n10059[4]; // extract
  assign n10443 = n10066[4]; // extract
  assign n10444 = n10071[4]; // extract
  assign n10445 = n10075[4]; // extract
  assign n10446 = n10078[4]; // extract
  assign n10447 = n10087[4]; // extract
  assign n10448 = n10179[4]; // extract
  assign n10449 = n10185[4]; // extract
  assign n10450 = n10217[4]; // extract
  assign n10451 = n10223[4]; // extract
  assign n10452 = n10255[4]; // extract
  assign n10453 = n10258[4]; // extract
  assign n10454 = n10261[4]; // extract
  assign n10455 = n10264[4]; // extract
  assign n10456 = n10267[4]; // extract
  assign n10457 = n10270[4]; // extract
  assign n10458 = n10273[4]; // extract
  assign n10459 = n10276[4]; // extract
  assign n10460 = n10279[4]; // extract
  assign n10461 = n10282[4]; // extract
  assign n10462 = n9998[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10463 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10463 = n10461;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10463 = n10460;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10463 = n10459;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10463 = n10458;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10463 = n10457;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10463 = n10456;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10463 = n10455;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10463 = n10454;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10463 = n10453;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10463 = n10452;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10463 = n10451;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10463 = n10450;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10463 = n10449;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10463 = n10448;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10463 = n10447;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10463 = n10446;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10463 = n10445;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10463 = n10444;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10463 = n10443;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10463 = n10442;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10463 = 1'b0;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10463 = n10441;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10463 = n10462;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10463 = n10462;
      default: n10463 = n10462;
    endcase
  assign n10464 = xcsr_rdata_i[5]; // extract
  assign n10465 = n10059[5]; // extract
  assign n10466 = n10066[5]; // extract
  assign n10467 = n10071[5]; // extract
  assign n10468 = n10078[5]; // extract
  assign n10469 = n10087[5]; // extract
  assign n10470 = n10179[5]; // extract
  assign n10471 = n10185[5]; // extract
  assign n10472 = n10217[5]; // extract
  assign n10473 = n10223[5]; // extract
  assign n10474 = n10255[5]; // extract
  assign n10475 = n10261[5]; // extract
  assign n10476 = n10264[5]; // extract
  assign n10477 = n10267[5]; // extract
  assign n10478 = n10270[5]; // extract
  assign n10479 = n10273[5]; // extract
  assign n10480 = n10276[5]; // extract
  assign n10481 = n10279[5]; // extract
  assign n10482 = n10282[5]; // extract
  assign n10483 = n9998[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10484 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10484 = n10482;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10484 = n10481;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10484 = n10480;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10484 = n10479;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10484 = n10478;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10484 = n10477;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10484 = n10476;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10484 = n10475;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10484 = n10474;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10484 = n10473;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10484 = n10472;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10484 = n10471;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10484 = n10470;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10484 = n10469;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10484 = n10468;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10484 = n10467;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10484 = n10466;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10484 = n10465;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10484 = n10464;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10484 = n10483;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10484 = n10483;
      default: n10484 = n10483;
    endcase
  assign n10485 = xcsr_rdata_i[6]; // extract
  assign n10486 = n10059[6]; // extract
  assign n10487 = n10066[6]; // extract
  assign n10488 = n10071[6]; // extract
  assign n10489 = n10078[6]; // extract
  assign n10490 = n10087[6]; // extract
  assign n10491 = n10179[6]; // extract
  assign n10492 = n10185[6]; // extract
  assign n10493 = n10217[6]; // extract
  assign n10494 = n10223[6]; // extract
  assign n10495 = n10255[6]; // extract
  assign n10496 = n10261[6]; // extract
  assign n10497 = n10264[6]; // extract
  assign n10498 = n10267[6]; // extract
  assign n10499 = n10270[6]; // extract
  assign n10500 = n10273[6]; // extract
  assign n10501 = n10276[6]; // extract
  assign n10502 = n10279[6]; // extract
  assign n10503 = n10282[6]; // extract
  assign n10504 = n9998[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10505 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10505 = n10503;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10505 = n10502;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10505 = n10501;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10505 = n10500;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10505 = n10499;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10505 = n10498;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10505 = n10497;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10505 = n10496;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10505 = n10495;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10505 = n10494;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10505 = n10493;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10505 = n10492;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10505 = n10491;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10505 = n10490;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10505 = n10489;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10505 = n10488;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10505 = n10487;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10505 = n10486;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10505 = n10485;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10505 = n10504;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10505 = n10504;
      default: n10505 = n10504;
    endcase
  assign n10506 = xcsr_rdata_i[7]; // extract
  assign n10507 = n10059[7]; // extract
  assign n10508 = n10066[7]; // extract
  assign n10509 = n10071[7]; // extract
  assign n10510 = n10078[7]; // extract
  assign n10511 = n10087[7]; // extract
  assign n10512 = n10179[7]; // extract
  assign n10513 = n10185[7]; // extract
  assign n10514 = n10217[7]; // extract
  assign n10515 = n10223[7]; // extract
  assign n10516 = n10255[7]; // extract
  assign n10517 = n10261[7]; // extract
  assign n10518 = n10264[7]; // extract
  assign n10519 = n10267[7]; // extract
  assign n10520 = n10270[7]; // extract
  assign n10521 = n10273[7]; // extract
  assign n10522 = n10276[7]; // extract
  assign n10523 = n10279[7]; // extract
  assign n10524 = n10282[7]; // extract
  assign n10525 = n9998[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10526 = 1'b1;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10526 = n10524;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10526 = n10523;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10526 = n10522;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10526 = n10521;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10526 = n10520;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10526 = n10519;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10526 = n10518;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10526 = n10517;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10526 = n10516;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10526 = n10515;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10526 = n10514;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10526 = n10513;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10526 = n10512;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10526 = n10511;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10526 = n10082;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10526 = n10510;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10526 = n10509;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10526 = n10508;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10526 = n10507;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10526 = n10054;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10526 = n10026;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10526 = n10506;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10526 = n10525;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10526 = n10525;
      default: n10526 = n10525;
    endcase
  assign n10527 = xcsr_rdata_i[8]; // extract
  assign n10528 = n10059[8]; // extract
  assign n10529 = n10066[8]; // extract
  assign n10530 = n10071[8]; // extract
  assign n10531 = n10078[8]; // extract
  assign n10532 = n10087[8]; // extract
  assign n10533 = n10179[8]; // extract
  assign n10534 = n10185[8]; // extract
  assign n10535 = n10217[8]; // extract
  assign n10536 = n10223[8]; // extract
  assign n10537 = n10255[8]; // extract
  assign n10538 = n10261[8]; // extract
  assign n10539 = n10264[8]; // extract
  assign n10540 = n10267[8]; // extract
  assign n10541 = n10270[8]; // extract
  assign n10542 = n10273[8]; // extract
  assign n10543 = n10276[8]; // extract
  assign n10544 = n10279[8]; // extract
  assign n10545 = n10282[8]; // extract
  assign n10546 = n9998[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10547 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10547 = n10545;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10547 = n10544;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10547 = n10543;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10547 = n10542;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10547 = n10541;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10547 = n10540;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10547 = n10539;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10547 = n10538;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10547 = n10537;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10547 = n10536;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10547 = n10535;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10547 = n10534;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10547 = n10533;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10547 = n10532;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10547 = n10531;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10547 = n10530;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10547 = n10529;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10547 = n10528;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10547 = 1'b1;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10547 = n10527;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10547 = n10546;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10547 = n10546;
      default: n10547 = n10546;
    endcase
  assign n10548 = xcsr_rdata_i[9]; // extract
  assign n10549 = n10059[9]; // extract
  assign n10550 = n10066[9]; // extract
  assign n10551 = n10071[9]; // extract
  assign n10552 = n10078[9]; // extract
  assign n10553 = n10087[9]; // extract
  assign n10554 = n10179[9]; // extract
  assign n10555 = n10185[9]; // extract
  assign n10556 = n10217[9]; // extract
  assign n10557 = n10223[9]; // extract
  assign n10558 = n10255[9]; // extract
  assign n10559 = n10261[9]; // extract
  assign n10560 = n10264[9]; // extract
  assign n10561 = n10267[9]; // extract
  assign n10562 = n10270[9]; // extract
  assign n10563 = n10273[9]; // extract
  assign n10564 = n10276[9]; // extract
  assign n10565 = n10279[9]; // extract
  assign n10566 = n10282[9]; // extract
  assign n10567 = n9998[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10568 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10568 = n10566;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10568 = n10565;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10568 = n10564;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10568 = n10563;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10568 = n10562;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10568 = n10561;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10568 = n10560;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10568 = n10559;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10568 = n10558;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10568 = n10557;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10568 = n10556;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10568 = n10555;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10568 = n10554;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10568 = n10553;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10568 = n10552;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10568 = n10551;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10568 = n10550;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10568 = n10549;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10568 = n10548;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10568 = n10567;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10568 = n10567;
      default: n10568 = n10567;
    endcase
  assign n10569 = xcsr_rdata_i[10]; // extract
  assign n10570 = n10059[10]; // extract
  assign n10571 = n10066[10]; // extract
  assign n10572 = n10071[10]; // extract
  assign n10573 = n10078[10]; // extract
  assign n10574 = n10087[10]; // extract
  assign n10575 = n10179[10]; // extract
  assign n10576 = n10185[10]; // extract
  assign n10577 = n10217[10]; // extract
  assign n10578 = n10223[10]; // extract
  assign n10579 = n10255[10]; // extract
  assign n10580 = n10261[10]; // extract
  assign n10581 = n10267[10]; // extract
  assign n10582 = n10270[10]; // extract
  assign n10583 = n10273[10]; // extract
  assign n10584 = n10276[10]; // extract
  assign n10585 = n10279[10]; // extract
  assign n10586 = n10282[10]; // extract
  assign n10587 = n9998[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10588 = 1'b1;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10588 = n10586;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10588 = n10585;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10588 = n10584;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10588 = n10583;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10588 = n10582;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10588 = n10581;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10588 = n10580;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10588 = n10579;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10588 = n10578;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10588 = n10577;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10588 = n10576;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10588 = n10575;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10588 = n10574;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10588 = n10573;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10588 = n10572;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10588 = n10571;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10588 = n10570;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10588 = n10569;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10588 = n10587;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10588 = n10587;
      default: n10588 = n10587;
    endcase
  assign n10589 = xcsr_rdata_i[11]; // extract
  assign n10590 = n10029[0]; // extract
  assign n10591 = n10059[11]; // extract
  assign n10592 = n10066[11]; // extract
  assign n10593 = n10071[11]; // extract
  assign n10594 = n10078[11]; // extract
  assign n10595 = n10087[11]; // extract
  assign n10596 = n10179[11]; // extract
  assign n10597 = n10185[11]; // extract
  assign n10598 = n10217[11]; // extract
  assign n10599 = n10223[11]; // extract
  assign n10600 = n10255[11]; // extract
  assign n10601 = n10261[11]; // extract
  assign n10602 = n10267[11]; // extract
  assign n10603 = n10270[11]; // extract
  assign n10604 = n10273[11]; // extract
  assign n10605 = n10276[11]; // extract
  assign n10606 = n10279[11]; // extract
  assign n10607 = n10282[11]; // extract
  assign n10608 = n9998[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10609 = 1'b1;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10609 = n10607;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10609 = n10606;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10609 = n10605;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10609 = n10604;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10609 = n10603;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10609 = n10602;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10609 = n10601;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10609 = n10600;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10609 = n10599;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10609 = n10598;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10609 = n10597;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10609 = n10596;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10609 = n10595;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10609 = n10083;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10609 = n10594;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10609 = n10593;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10609 = n10592;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10609 = n10591;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10609 = n10055;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10609 = n10590;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10609 = n10589;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10609 = n10608;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10609 = n10608;
      default: n10609 = n10608;
    endcase
  assign n10610 = xcsr_rdata_i[12]; // extract
  assign n10611 = n10029[1]; // extract
  assign n10612 = n10059[12]; // extract
  assign n10613 = n10066[12]; // extract
  assign n10614 = n10071[12]; // extract
  assign n10615 = n10078[12]; // extract
  assign n10616 = n10087[12]; // extract
  assign n10617 = n10179[12]; // extract
  assign n10618 = n10185[12]; // extract
  assign n10619 = n10217[12]; // extract
  assign n10620 = n10223[12]; // extract
  assign n10621 = n10255[12]; // extract
  assign n10622 = n10261[12]; // extract
  assign n10623 = n10267[12]; // extract
  assign n10624 = n10270[12]; // extract
  assign n10625 = n10273[12]; // extract
  assign n10626 = n10276[12]; // extract
  assign n10627 = n10279[12]; // extract
  assign n10628 = n10282[12]; // extract
  assign n10629 = n9998[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10630 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10630 = n10628;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10630 = n10627;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10630 = n10626;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10630 = n10625;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10630 = n10624;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10630 = n10623;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10630 = n10622;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10630 = n10621;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10630 = n10620;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10630 = n10619;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10630 = n10618;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10630 = n10617;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10630 = n10616;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10630 = n10615;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10630 = n10614;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10630 = n10613;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10630 = n10612;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10630 = 1'b1;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10630 = n10611;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10630 = n10610;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10630 = n10629;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10630 = n10629;
      default: n10630 = n10629;
    endcase
  assign n10631 = xcsr_rdata_i[13]; // extract
  assign n10632 = n10059[13]; // extract
  assign n10633 = n10066[13]; // extract
  assign n10634 = n10071[13]; // extract
  assign n10635 = n10078[13]; // extract
  assign n10636 = n10087[13]; // extract
  assign n10637 = n10179[13]; // extract
  assign n10638 = n10185[13]; // extract
  assign n10639 = n10217[13]; // extract
  assign n10640 = n10223[13]; // extract
  assign n10641 = n10255[13]; // extract
  assign n10642 = n10261[13]; // extract
  assign n10643 = n10267[13]; // extract
  assign n10644 = n10270[13]; // extract
  assign n10645 = n10273[13]; // extract
  assign n10646 = n10276[13]; // extract
  assign n10647 = n10279[13]; // extract
  assign n10648 = n10282[13]; // extract
  assign n10649 = n9998[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10650 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10650 = n10648;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10650 = n10647;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10650 = n10646;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10650 = n10645;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10650 = n10644;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10650 = n10643;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10650 = n10642;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10650 = n10641;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10650 = n10640;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10650 = n10639;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10650 = n10638;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10650 = n10637;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10650 = n10636;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10650 = n10635;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10650 = n10634;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10650 = n10633;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10650 = n10632;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10650 = n10631;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10650 = n10649;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10650 = n10649;
      default: n10650 = n10649;
    endcase
  assign n10651 = xcsr_rdata_i[14]; // extract
  assign n10652 = n10059[14]; // extract
  assign n10653 = n10066[14]; // extract
  assign n10654 = n10071[14]; // extract
  assign n10655 = n10078[14]; // extract
  assign n10656 = n10087[14]; // extract
  assign n10657 = n10179[14]; // extract
  assign n10658 = n10185[14]; // extract
  assign n10659 = n10217[14]; // extract
  assign n10660 = n10223[14]; // extract
  assign n10661 = n10255[14]; // extract
  assign n10662 = n10261[14]; // extract
  assign n10663 = n10267[14]; // extract
  assign n10664 = n10270[14]; // extract
  assign n10665 = n10273[14]; // extract
  assign n10666 = n10276[14]; // extract
  assign n10667 = n10279[14]; // extract
  assign n10668 = n10282[14]; // extract
  assign n10669 = n9998[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10670 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10670 = n10668;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10670 = n10667;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10670 = n10666;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10670 = n10665;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10670 = n10664;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10670 = n10663;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10670 = n10662;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10670 = n10661;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10670 = n10660;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10670 = n10659;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10670 = n10658;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10670 = n10657;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10670 = n10656;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10670 = n10655;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10670 = n10654;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10670 = n10653;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10670 = n10652;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10670 = n10651;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10670 = n10669;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10670 = n10669;
      default: n10670 = n10669;
    endcase
  assign n10671 = xcsr_rdata_i[15]; // extract
  assign n10672 = n10059[15]; // extract
  assign n10673 = n10066[15]; // extract
  assign n10674 = n10071[15]; // extract
  assign n10675 = n10078[15]; // extract
  assign n10676 = n10087[15]; // extract
  assign n10677 = n10179[15]; // extract
  assign n10678 = n10185[15]; // extract
  assign n10679 = n10217[15]; // extract
  assign n10680 = n10223[15]; // extract
  assign n10681 = n10255[15]; // extract
  assign n10682 = n10261[15]; // extract
  assign n10683 = n10267[15]; // extract
  assign n10684 = n10270[15]; // extract
  assign n10685 = n10273[15]; // extract
  assign n10686 = n10276[15]; // extract
  assign n10687 = n10279[15]; // extract
  assign n10688 = n10282[15]; // extract
  assign n10689 = n9998[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10690 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10690 = n10688;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10690 = n10687;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10690 = n10686;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10690 = n10685;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10690 = n10684;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10690 = n10683;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10690 = n10682;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10690 = n10681;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10690 = n10680;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10690 = n10679;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10690 = n10678;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10690 = n10677;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10690 = n10676;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10690 = n10675;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10690 = n10674;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10690 = n10673;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10690 = n10672;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10690 = n10671;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10690 = n10689;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10690 = n10689;
      default: n10690 = n10689;
    endcase
  assign n10691 = xcsr_rdata_i[16]; // extract
  assign n10692 = n10056[0]; // extract
  assign n10693 = n10059[16]; // extract
  assign n10694 = n10066[16]; // extract
  assign n10695 = n10071[16]; // extract
  assign n10696 = n10078[16]; // extract
  assign n10697 = n10084[0]; // extract
  assign n10698 = n10087[16]; // extract
  assign n10699 = n10179[16]; // extract
  assign n10700 = n10185[16]; // extract
  assign n10701 = n10217[16]; // extract
  assign n10702 = n10223[16]; // extract
  assign n10703 = n10255[16]; // extract
  assign n10704 = n10261[16]; // extract
  assign n10705 = n10267[16]; // extract
  assign n10706 = n10270[16]; // extract
  assign n10707 = n10273[16]; // extract
  assign n10708 = n10276[16]; // extract
  assign n10709 = n10279[16]; // extract
  assign n10710 = n10282[16]; // extract
  assign n10711 = n9998[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10712 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10712 = n10710;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10712 = n10709;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10712 = n10708;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10712 = n10707;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10712 = n10706;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10712 = n10705;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10712 = n10704;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10712 = n10703;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10712 = n10702;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10712 = n10701;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10712 = n10700;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10712 = n10699;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10712 = n10698;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10712 = n10697;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10712 = n10696;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10712 = n10695;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10712 = n10694;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10712 = n10693;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10712 = n10692;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10712 = n10691;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10712 = n10711;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10712 = n10711;
      default: n10712 = n10711;
    endcase
  assign n10713 = xcsr_rdata_i[17]; // extract
  assign n10714 = n10056[1]; // extract
  assign n10715 = n10059[17]; // extract
  assign n10716 = n10066[17]; // extract
  assign n10717 = n10071[17]; // extract
  assign n10718 = n10078[17]; // extract
  assign n10719 = n10084[1]; // extract
  assign n10720 = n10087[17]; // extract
  assign n10721 = n10179[17]; // extract
  assign n10722 = n10185[17]; // extract
  assign n10723 = n10217[17]; // extract
  assign n10724 = n10223[17]; // extract
  assign n10725 = n10255[17]; // extract
  assign n10726 = n10261[17]; // extract
  assign n10727 = n10267[17]; // extract
  assign n10728 = n10270[17]; // extract
  assign n10729 = n10273[17]; // extract
  assign n10730 = n10276[17]; // extract
  assign n10731 = n10279[17]; // extract
  assign n10732 = n10282[17]; // extract
  assign n10733 = n9998[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10734 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10734 = n10732;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10734 = n10731;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10734 = n10730;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10734 = n10729;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10734 = n10728;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10734 = n10727;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10734 = n10726;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10734 = n10725;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10734 = n10724;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10734 = n10723;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10734 = n10722;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10734 = n10721;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10734 = n10720;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10734 = n10719;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10734 = n10718;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10734 = n10717;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10734 = n10716;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10734 = n10715;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10734 = n10714;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10734 = n10030;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10734 = n10713;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10734 = n10733;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10734 = n10733;
      default: n10734 = n10733;
    endcase
  assign n10735 = xcsr_rdata_i[18]; // extract
  assign n10736 = n10056[2]; // extract
  assign n10737 = n10059[18]; // extract
  assign n10738 = n10066[18]; // extract
  assign n10739 = n10071[18]; // extract
  assign n10740 = n10078[18]; // extract
  assign n10741 = n10084[2]; // extract
  assign n10742 = n10087[18]; // extract
  assign n10743 = n10179[18]; // extract
  assign n10744 = n10185[18]; // extract
  assign n10745 = n10217[18]; // extract
  assign n10746 = n10223[18]; // extract
  assign n10747 = n10255[18]; // extract
  assign n10748 = n10261[18]; // extract
  assign n10749 = n10267[18]; // extract
  assign n10750 = n10270[18]; // extract
  assign n10751 = n10273[18]; // extract
  assign n10752 = n10276[18]; // extract
  assign n10753 = n10279[18]; // extract
  assign n10754 = n10282[18]; // extract
  assign n10755 = n9998[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10756 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10756 = n10754;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10756 = n10753;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10756 = n10752;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10756 = n10751;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10756 = n10750;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10756 = n10749;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10756 = n10748;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10756 = n10747;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10756 = n10746;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10756 = n10745;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10756 = n10744;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10756 = n10743;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10756 = n10742;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10756 = n10741;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10756 = n10740;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10756 = n10739;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10756 = n10738;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10756 = n10737;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10756 = n10736;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10756 = n10735;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10756 = n10755;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10756 = n10755;
      default: n10756 = n10755;
    endcase
  assign n10757 = xcsr_rdata_i[19]; // extract
  assign n10758 = n10056[3]; // extract
  assign n10759 = n10059[19]; // extract
  assign n10760 = n10066[19]; // extract
  assign n10761 = n10071[19]; // extract
  assign n10762 = n10078[19]; // extract
  assign n10763 = n10084[3]; // extract
  assign n10764 = n10087[19]; // extract
  assign n10765 = n10179[19]; // extract
  assign n10766 = n10185[19]; // extract
  assign n10767 = n10217[19]; // extract
  assign n10768 = n10223[19]; // extract
  assign n10769 = n10255[19]; // extract
  assign n10770 = n10261[19]; // extract
  assign n10771 = n10267[19]; // extract
  assign n10772 = n10270[19]; // extract
  assign n10773 = n10273[19]; // extract
  assign n10774 = n10276[19]; // extract
  assign n10775 = n10279[19]; // extract
  assign n10776 = n10282[19]; // extract
  assign n10777 = n9998[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10778 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10778 = n10776;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10778 = n10775;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10778 = n10774;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10778 = n10773;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10778 = n10772;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10778 = n10771;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10778 = n10770;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10778 = n10769;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10778 = n10768;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10778 = n10767;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10778 = n10766;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10778 = n10765;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10778 = n10764;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10778 = n10763;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10778 = n10762;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10778 = n10761;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10778 = n10760;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10778 = n10759;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10778 = n10758;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10778 = n10757;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10778 = n10777;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10778 = n10777;
      default: n10778 = n10777;
    endcase
  assign n10779 = xcsr_rdata_i[20]; // extract
  assign n10780 = n10056[4]; // extract
  assign n10781 = n10059[20]; // extract
  assign n10782 = n10066[20]; // extract
  assign n10783 = n10071[20]; // extract
  assign n10784 = n10078[20]; // extract
  assign n10785 = n10084[4]; // extract
  assign n10786 = n10087[20]; // extract
  assign n10787 = n10179[20]; // extract
  assign n10788 = n10185[20]; // extract
  assign n10789 = n10217[20]; // extract
  assign n10790 = n10223[20]; // extract
  assign n10791 = n10255[20]; // extract
  assign n10792 = n10261[20]; // extract
  assign n10793 = n10267[20]; // extract
  assign n10794 = n10270[20]; // extract
  assign n10795 = n10273[20]; // extract
  assign n10796 = n10276[20]; // extract
  assign n10797 = n10279[20]; // extract
  assign n10798 = n10282[20]; // extract
  assign n10799 = n9998[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10800 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10800 = n10798;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10800 = n10797;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10800 = n10796;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10800 = n10795;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10800 = n10794;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10800 = n10793;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10800 = n10792;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10800 = n10791;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10800 = n10790;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10800 = n10789;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10800 = n10788;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10800 = n10787;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10800 = n10786;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10800 = n10785;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10800 = n10784;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10800 = n10783;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10800 = n10782;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10800 = n10781;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10800 = n10780;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10800 = 1'b1;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10800 = n10779;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10800 = n10799;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10800 = n10799;
      default: n10800 = n10799;
    endcase
  assign n10801 = xcsr_rdata_i[21]; // extract
  assign n10802 = n10056[5]; // extract
  assign n10803 = n10059[21]; // extract
  assign n10804 = n10066[21]; // extract
  assign n10805 = n10071[21]; // extract
  assign n10806 = n10078[21]; // extract
  assign n10807 = n10084[5]; // extract
  assign n10808 = n10087[21]; // extract
  assign n10809 = n10179[21]; // extract
  assign n10810 = n10185[21]; // extract
  assign n10811 = n10217[21]; // extract
  assign n10812 = n10223[21]; // extract
  assign n10813 = n10255[21]; // extract
  assign n10814 = n10261[21]; // extract
  assign n10815 = n10267[21]; // extract
  assign n10816 = n10270[21]; // extract
  assign n10817 = n10273[21]; // extract
  assign n10818 = n10276[21]; // extract
  assign n10819 = n10279[21]; // extract
  assign n10820 = n10282[21]; // extract
  assign n10821 = n9998[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10822 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10822 = n10820;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10822 = n10819;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10822 = n10818;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10822 = n10817;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10822 = n10816;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10822 = n10815;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10822 = n10814;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10822 = n10813;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10822 = n10812;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10822 = n10811;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10822 = n10810;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10822 = n10809;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10822 = n10808;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10822 = n10807;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10822 = n10806;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10822 = n10805;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10822 = n10804;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10822 = n10803;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10822 = n10802;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10822 = n10034;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10822 = n10801;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10822 = n10821;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10822 = n10821;
      default: n10822 = n10821;
    endcase
  assign n10823 = xcsr_rdata_i[22]; // extract
  assign n10824 = n10056[6]; // extract
  assign n10825 = n10059[22]; // extract
  assign n10826 = n10066[22]; // extract
  assign n10827 = n10071[22]; // extract
  assign n10828 = n10078[22]; // extract
  assign n10829 = n10084[6]; // extract
  assign n10830 = n10087[22]; // extract
  assign n10831 = n10179[22]; // extract
  assign n10832 = n10185[22]; // extract
  assign n10833 = n10217[22]; // extract
  assign n10834 = n10223[22]; // extract
  assign n10835 = n10255[22]; // extract
  assign n10836 = n10261[22]; // extract
  assign n10837 = n10267[22]; // extract
  assign n10838 = n10270[22]; // extract
  assign n10839 = n10273[22]; // extract
  assign n10840 = n10276[22]; // extract
  assign n10841 = n10279[22]; // extract
  assign n10842 = n10282[22]; // extract
  assign n10843 = n9998[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10844 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10844 = n10842;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10844 = n10841;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10844 = n10840;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10844 = n10839;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10844 = n10838;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10844 = n10837;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10844 = n10836;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10844 = n10835;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10844 = n10834;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10844 = n10833;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10844 = n10832;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10844 = n10831;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10844 = n10830;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10844 = n10829;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10844 = n10828;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10844 = n10827;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10844 = n10826;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10844 = n10825;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10844 = n10824;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10844 = n10823;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10844 = n10843;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10844 = n10843;
      default: n10844 = n10843;
    endcase
  assign n10845 = xcsr_rdata_i[23]; // extract
  assign n10846 = n10056[7]; // extract
  assign n10847 = n10059[23]; // extract
  assign n10848 = n10066[23]; // extract
  assign n10849 = n10071[23]; // extract
  assign n10850 = n10078[23]; // extract
  assign n10851 = n10084[7]; // extract
  assign n10852 = n10087[23]; // extract
  assign n10853 = n10179[23]; // extract
  assign n10854 = n10185[23]; // extract
  assign n10855 = n10217[23]; // extract
  assign n10856 = n10223[23]; // extract
  assign n10857 = n10255[23]; // extract
  assign n10858 = n10261[23]; // extract
  assign n10859 = n10267[23]; // extract
  assign n10860 = n10270[23]; // extract
  assign n10861 = n10273[23]; // extract
  assign n10862 = n10276[23]; // extract
  assign n10863 = n10279[23]; // extract
  assign n10864 = n10282[23]; // extract
  assign n10865 = n9998[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10866 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10866 = n10864;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10866 = n10863;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10866 = n10862;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10866 = n10861;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10866 = n10860;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10866 = n10859;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10866 = n10858;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10866 = n10857;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10866 = n10856;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10866 = n10855;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10866 = n10854;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10866 = n10853;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10866 = n10852;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10866 = n10851;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10866 = n10850;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10866 = n10849;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10866 = n10848;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10866 = n10847;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10866 = n10846;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10866 = 1'b1;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10866 = n10845;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10866 = n10865;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10866 = n10865;
      default: n10866 = n10865;
    endcase
  assign n10867 = xcsr_rdata_i[24]; // extract
  assign n10868 = n10056[8]; // extract
  assign n10869 = n10059[24]; // extract
  assign n10870 = n10066[24]; // extract
  assign n10871 = n10071[24]; // extract
  assign n10872 = n10078[24]; // extract
  assign n10873 = n10084[8]; // extract
  assign n10874 = n10087[24]; // extract
  assign n10875 = n10179[24]; // extract
  assign n10876 = n10185[24]; // extract
  assign n10877 = n10217[24]; // extract
  assign n10878 = n10223[24]; // extract
  assign n10879 = n10255[24]; // extract
  assign n10880 = n10261[24]; // extract
  assign n10881 = n10267[24]; // extract
  assign n10882 = n10270[24]; // extract
  assign n10883 = n10273[24]; // extract
  assign n10884 = n10276[24]; // extract
  assign n10885 = n10279[24]; // extract
  assign n10886 = n10282[24]; // extract
  assign n10887 = n9998[24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10888 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10888 = n10886;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10888 = n10885;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10888 = n10884;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10888 = n10883;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10888 = n10882;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10888 = n10881;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10888 = n10880;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10888 = n10879;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10888 = n10878;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10888 = n10877;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10888 = n10876;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10888 = n10875;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10888 = n10874;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10888 = n10873;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10888 = n10872;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10888 = n10871;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10888 = n10870;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10888 = n10869;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10888 = n10868;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10888 = n10867;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10888 = n10887;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10888 = n10887;
      default: n10888 = n10887;
    endcase
  assign n10889 = xcsr_rdata_i[25]; // extract
  assign n10890 = n10056[9]; // extract
  assign n10891 = n10059[25]; // extract
  assign n10892 = n10066[25]; // extract
  assign n10893 = n10071[25]; // extract
  assign n10894 = n10078[25]; // extract
  assign n10895 = n10084[9]; // extract
  assign n10896 = n10087[25]; // extract
  assign n10897 = n10179[25]; // extract
  assign n10898 = n10185[25]; // extract
  assign n10899 = n10217[25]; // extract
  assign n10900 = n10223[25]; // extract
  assign n10901 = n10255[25]; // extract
  assign n10902 = n10261[25]; // extract
  assign n10903 = n10267[25]; // extract
  assign n10904 = n10270[25]; // extract
  assign n10905 = n10273[25]; // extract
  assign n10906 = n10276[25]; // extract
  assign n10907 = n10279[25]; // extract
  assign n10908 = n10282[25]; // extract
  assign n10909 = n9998[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10910 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10910 = n10908;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10910 = n10907;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10910 = n10906;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10910 = n10905;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10910 = n10904;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10910 = n10903;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10910 = n10902;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10910 = n10901;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10910 = n10900;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10910 = n10899;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10910 = n10898;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10910 = n10897;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10910 = n10896;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10910 = n10895;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10910 = n10894;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10910 = n10893;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10910 = n10892;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10910 = n10891;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10910 = n10890;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10910 = n10889;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10910 = n10909;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10910 = n10909;
      default: n10910 = n10909;
    endcase
  assign n10911 = xcsr_rdata_i[26]; // extract
  assign n10912 = n10056[10]; // extract
  assign n10913 = n10059[26]; // extract
  assign n10914 = n10066[26]; // extract
  assign n10915 = n10071[26]; // extract
  assign n10916 = n10078[26]; // extract
  assign n10917 = n10084[10]; // extract
  assign n10918 = n10087[26]; // extract
  assign n10919 = n10179[26]; // extract
  assign n10920 = n10185[26]; // extract
  assign n10921 = n10217[26]; // extract
  assign n10922 = n10223[26]; // extract
  assign n10923 = n10255[26]; // extract
  assign n10924 = n10261[26]; // extract
  assign n10925 = n10267[26]; // extract
  assign n10926 = n10270[26]; // extract
  assign n10927 = n10273[26]; // extract
  assign n10928 = n10276[26]; // extract
  assign n10929 = n10279[26]; // extract
  assign n10930 = n10282[26]; // extract
  assign n10931 = n9998[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10932 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10932 = n10930;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10932 = n10929;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10932 = n10928;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10932 = n10927;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10932 = n10926;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10932 = n10925;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10932 = n10924;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10932 = n10923;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10932 = n10922;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10932 = n10921;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10932 = n10920;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10932 = n10919;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10932 = n10918;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10932 = n10917;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10932 = n10916;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10932 = n10915;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10932 = n10914;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10932 = n10913;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10932 = n10912;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10932 = n10911;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10932 = n10931;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10932 = n10931;
      default: n10932 = n10931;
    endcase
  assign n10933 = xcsr_rdata_i[27]; // extract
  assign n10934 = n10056[11]; // extract
  assign n10935 = n10059[27]; // extract
  assign n10936 = n10066[27]; // extract
  assign n10937 = n10071[27]; // extract
  assign n10938 = n10078[27]; // extract
  assign n10939 = n10084[11]; // extract
  assign n10940 = n10087[27]; // extract
  assign n10941 = n10179[27]; // extract
  assign n10942 = n10185[27]; // extract
  assign n10943 = n10217[27]; // extract
  assign n10944 = n10223[27]; // extract
  assign n10945 = n10255[27]; // extract
  assign n10946 = n10261[27]; // extract
  assign n10947 = n10267[27]; // extract
  assign n10948 = n10270[27]; // extract
  assign n10949 = n10273[27]; // extract
  assign n10950 = n10276[27]; // extract
  assign n10951 = n10279[27]; // extract
  assign n10952 = n10282[27]; // extract
  assign n10953 = n9998[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10954 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10954 = n10952;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10954 = n10951;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10954 = n10950;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10954 = n10949;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10954 = n10948;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10954 = n10947;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10954 = n10946;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10954 = n10945;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10954 = n10944;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10954 = n10943;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10954 = n10942;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10954 = n10941;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10954 = n10940;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10954 = n10939;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10954 = n10938;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10954 = n10937;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10954 = n10936;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10954 = n10935;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10954 = n10934;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10954 = n10933;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10954 = n10953;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10954 = n10953;
      default: n10954 = n10953;
    endcase
  assign n10955 = xcsr_rdata_i[28]; // extract
  assign n10956 = n10056[12]; // extract
  assign n10957 = n10059[28]; // extract
  assign n10958 = n10066[28]; // extract
  assign n10959 = n10071[28]; // extract
  assign n10960 = n10078[28]; // extract
  assign n10961 = n10084[12]; // extract
  assign n10962 = n10087[28]; // extract
  assign n10963 = n10179[28]; // extract
  assign n10964 = n10185[28]; // extract
  assign n10965 = n10217[28]; // extract
  assign n10966 = n10223[28]; // extract
  assign n10967 = n10255[28]; // extract
  assign n10968 = n10261[28]; // extract
  assign n10969 = n10267[28]; // extract
  assign n10970 = n10270[28]; // extract
  assign n10971 = n10273[28]; // extract
  assign n10972 = n10276[28]; // extract
  assign n10973 = n10279[28]; // extract
  assign n10974 = n10282[28]; // extract
  assign n10975 = n9998[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10976 = 1'b1;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10976 = n10974;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10976 = n10973;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10976 = n10972;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10976 = n10971;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10976 = n10970;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10976 = n10969;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10976 = n10968;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10976 = n10967;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10976 = n10966;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10976 = n10965;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10976 = n10964;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10976 = n10963;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10976 = n10962;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10976 = n10961;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10976 = n10960;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10976 = n10959;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10976 = n10958;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10976 = n10957;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10976 = n10956;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10976 = n10955;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10976 = n10975;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10976 = n10975;
      default: n10976 = n10975;
    endcase
  assign n10977 = xcsr_rdata_i[29]; // extract
  assign n10978 = n10056[13]; // extract
  assign n10979 = n10059[29]; // extract
  assign n10980 = n10066[29]; // extract
  assign n10981 = n10071[29]; // extract
  assign n10982 = n10078[29]; // extract
  assign n10983 = n10084[13]; // extract
  assign n10984 = n10087[29]; // extract
  assign n10985 = n10179[29]; // extract
  assign n10986 = n10185[29]; // extract
  assign n10987 = n10217[29]; // extract
  assign n10988 = n10223[29]; // extract
  assign n10989 = n10255[29]; // extract
  assign n10990 = n10261[29]; // extract
  assign n10991 = n10267[29]; // extract
  assign n10992 = n10270[29]; // extract
  assign n10993 = n10273[29]; // extract
  assign n10994 = n10276[29]; // extract
  assign n10995 = n10279[29]; // extract
  assign n10996 = n10282[29]; // extract
  assign n10997 = n9998[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n10998 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n10998 = n10996;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n10998 = n10995;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n10998 = n10994;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n10998 = n10993;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n10998 = n10992;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n10998 = n10991;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n10998 = n10990;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n10998 = n10989;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n10998 = n10988;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n10998 = n10987;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n10998 = n10986;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n10998 = n10985;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n10998 = n10984;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n10998 = n10983;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n10998 = n10982;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n10998 = n10981;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n10998 = n10980;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n10998 = n10979;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n10998 = n10978;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n10998 = n10977;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n10998 = n10997;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n10998 = n10997;
      default: n10998 = n10997;
    endcase
  assign n10999 = xcsr_rdata_i[30]; // extract
  assign n11000 = n10050[0]; // extract
  assign n11001 = n10056[14]; // extract
  assign n11002 = n10059[30]; // extract
  assign n11003 = n10066[30]; // extract
  assign n11004 = n10071[30]; // extract
  assign n11005 = n10078[30]; // extract
  assign n11006 = n10084[14]; // extract
  assign n11007 = n10087[30]; // extract
  assign n11008 = n10179[30]; // extract
  assign n11009 = n10185[30]; // extract
  assign n11010 = n10217[30]; // extract
  assign n11011 = n10223[30]; // extract
  assign n11012 = n10255[30]; // extract
  assign n11013 = n10261[30]; // extract
  assign n11014 = n10267[30]; // extract
  assign n11015 = n10270[30]; // extract
  assign n11016 = n10273[30]; // extract
  assign n11017 = n10276[30]; // extract
  assign n11018 = n10279[30]; // extract
  assign n11019 = n10282[30]; // extract
  assign n11020 = n9998[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n11021 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n11021 = n11019;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n11021 = n11018;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n11021 = n11017;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n11021 = n11016;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n11021 = n11015;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n11021 = n11014;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n11021 = n11013;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n11021 = n11012;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n11021 = n11011;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n11021 = n11010;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n11021 = n11009;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n11021 = n11008;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n11021 = n11007;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n11021 = n11006;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n11021 = n11005;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n11021 = n11004;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n11021 = n11003;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n11021 = n11002;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n11021 = n11001;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n11021 = n11000;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n11021 = n10999;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n11021 = n11020;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n11021 = n11020;
      default: n11021 = n11020;
    endcase
  assign n11022 = xcsr_rdata_i[31]; // extract
  assign n11023 = n10050[1]; // extract
  assign n11024 = n10056[15]; // extract
  assign n11025 = n10059[31]; // extract
  assign n11026 = n10066[31]; // extract
  assign n11027 = n10071[31]; // extract
  assign n11028 = n10078[31]; // extract
  assign n11029 = n10084[15]; // extract
  assign n11030 = n10087[31]; // extract
  assign n11031 = n10179[31]; // extract
  assign n11032 = n10185[31]; // extract
  assign n11033 = n10217[31]; // extract
  assign n11034 = n10223[31]; // extract
  assign n11035 = n10255[31]; // extract
  assign n11036 = n10261[31]; // extract
  assign n11037 = n10267[31]; // extract
  assign n11038 = n10270[31]; // extract
  assign n11039 = n10273[31]; // extract
  assign n11040 = n10276[31]; // extract
  assign n11041 = n10279[31]; // extract
  assign n11042 = n10282[31]; // extract
  assign n11043 = n9998[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1654:9  */
  always @*
    case (n10348)
      70'b1000000000000000000000000000000000000000000000000000000000000000000000: n11044 = 1'b0;
      70'b0100000000000000000000000000000000000000000000000000000000000000000000: n11044 = n11042;
      70'b0010000000000000000000000000000000000000000000000000000000000000000000: n11044 = n11041;
      70'b0001000000000000000000000000000000000000000000000000000000000000000000: n11044 = n11040;
      70'b0000100000000000000000000000000000000000000000000000000000000000000000: n11044 = n11039;
      70'b0000010000000000000000000000000000000000000000000000000000000000000000: n11044 = n11038;
      70'b0000001000000000000000000000000000000000000000000000000000000000000000: n11044 = n11037;
      70'b0000000100000000000000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000010000000000000000000000000000000000000000000000000000000000000: n11044 = n11036;
      70'b0000000001000000000000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000100000000000000000000000000000000000000000000000000000000000: n11044 = n11035;
      70'b0000000000010000000000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000001000000000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000100000000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000010000000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000001000000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000100000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000010000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000001000000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000100000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000010000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000001000000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000100000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000010000000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000001000000000000000000000000000000000000000000000: n11044 = n11034;
      70'b0000000000000000000000000100000000000000000000000000000000000000000000: n11044 = n11033;
      70'b0000000000000000000000000010000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000001000000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000100000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000010000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000001000000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000100000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000010000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000001000000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000100000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000010000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000001000000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000100000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000010000000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000001000000000000000000000000000000: n11044 = n11032;
      70'b0000000000000000000000000000000000000000100000000000000000000000000000: n11044 = n11031;
      70'b0000000000000000000000000000000000000000010000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000001000000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000100000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000010000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000001000000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000100000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000010000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000001000000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000100000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000010000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000001000000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000000100000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000000010000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000000001000000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000000000100000000000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000000000010000000000000: n11044 = n11030;
      70'b0000000000000000000000000000000000000000000000000000000001000000000000: n11044 = n11029;
      70'b0000000000000000000000000000000000000000000000000000000000100000000000: n11044 = n11028;
      70'b0000000000000000000000000000000000000000000000000000000000010000000000: n11044 = n10074;
      70'b0000000000000000000000000000000000000000000000000000000000001000000000: n11044 = n11027;
      70'b0000000000000000000000000000000000000000000000000000000000000100000000: n11044 = n11026;
      70'b0000000000000000000000000000000000000000000000000000000000000010000000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000000000000000001000000: n11044 = n11025;
      70'b0000000000000000000000000000000000000000000000000000000000000000100000: n11044 = n11024;
      70'b0000000000000000000000000000000000000000000000000000000000000000010000: n11044 = n11023;
      70'b0000000000000000000000000000000000000000000000000000000000000000001000: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000000000000000000000100: n11044 = n11022;
      70'b0000000000000000000000000000000000000000000000000000000000000000000010: n11044 = n11043;
      70'b0000000000000000000000000000000000000000000000000000000000000000000001: n11044 = n11043;
      default: n11044 = n11043;
    endcase
  assign n11045 = {n11044, n11021, n10998, n10976, n10954, n10932, n10910, n10888, n10866, n10844, n10822, n10800, n10778, n10756, n10734, n10712, n10690, n10670, n10650, n10630, n10609, n10588, n10568, n10547, n10526, n10505, n10484, n10463, n10440, n10417, n10394, n10371};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1653:7  */
  assign n11046 = n9999 ? n11045 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1900:22  */
  assign n11054 = csr[111:80]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:18  */
  assign n11056 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:17  */
  assign n11061 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:40  */
  assign n11062 = csr[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:54  */
  assign n11064 = n11062 == 5'b10110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:27  */
  assign n11065 = n11064 & n11061;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1923:21  */
  assign n11066 = csr[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1923:34  */
  assign n11068 = n11066 == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:83  */
  assign n11069 = n11068 & n11065;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1924:28  */
  assign n11070 = csr[79:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1926:34  */
  assign n11071 = cnt[305:274]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:9  */
  assign n11072 = n11069 ? n11070 : n11071;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1928:36  */
  assign n11073 = cnt[306]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:17  */
  assign n11074 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:40  */
  assign n11075 = csr[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:54  */
  assign n11077 = n11075 == 5'b10111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:27  */
  assign n11078 = n11077 & n11074;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1932:21  */
  assign n11079 = csr[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1932:34  */
  assign n11081 = n11079 == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:84  */
  assign n11082 = n11081 & n11078;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1933:28  */
  assign n11083 = csr[79:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:57  */
  assign n11084 = cnt[207:176]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:80  */
  assign n11085 = cnt[309]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:62  */
  assign n11086 = {31'b0, n11085};  //  uext
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:62  */
  assign n11087 = n11084 + n11086;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:9  */
  assign n11088 = n11082 ? n11083 : n11087;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:58  */
  assign n11099 = cnt[111:80]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:50  */
  assign n11101 = {1'b0, n11099};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:81  */
  assign n11102 = cnt[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:63  */
  assign n11103 = {32'b0, n11102};  //  uext
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:63  */
  assign n11104 = n11101 + n11103;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:18  */
  assign n11106 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:17  */
  assign n11111 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:40  */
  assign n11112 = csr[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:54  */
  assign n11114 = n11112 == 5'b10110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:27  */
  assign n11115 = n11114 & n11111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1923:21  */
  assign n11116 = csr[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1923:34  */
  assign n11118 = n11116 == 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:83  */
  assign n11119 = n11118 & n11115;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1924:28  */
  assign n11120 = csr[79:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1926:34  */
  assign n11121 = cnt[272:241]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:9  */
  assign n11122 = n11119 ? n11120 : n11121;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1928:36  */
  assign n11123 = cnt[273]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:17  */
  assign n11124 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:40  */
  assign n11125 = csr[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:54  */
  assign n11127 = n11125 == 5'b10111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:27  */
  assign n11128 = n11127 & n11124;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1932:21  */
  assign n11129 = csr[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1932:34  */
  assign n11131 = n11129 == 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:84  */
  assign n11132 = n11131 & n11128;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1933:28  */
  assign n11133 = csr[79:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:57  */
  assign n11134 = cnt[175:144]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:80  */
  assign n11135 = cnt[308]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:62  */
  assign n11136 = {31'b0, n11135};  //  uext
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:62  */
  assign n11137 = n11134 + n11136;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:9  */
  assign n11138 = n11132 ? n11133 : n11137;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:58  */
  assign n11149 = cnt[79:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:50  */
  assign n11151 = {1'b0, n11149};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:81  */
  assign n11152 = cnt[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:63  */
  assign n11153 = {32'b0, n11152};  //  uext
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:63  */
  assign n11154 = n11151 + n11153;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:18  */
  assign n11156 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:17  */
  assign n11161 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:40  */
  assign n11162 = csr[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:54  */
  assign n11164 = n11162 == 5'b10110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:27  */
  assign n11165 = n11164 & n11161;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1923:21  */
  assign n11166 = csr[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1923:34  */
  assign n11168 = n11166 == 4'b0010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:83  */
  assign n11169 = n11168 & n11165;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1924:28  */
  assign n11170 = csr[79:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1926:34  */
  assign n11171 = cnt[239:208]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1922:9  */
  assign n11172 = n11169 ? n11170 : n11171;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1928:36  */
  assign n11173 = cnt[240]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:17  */
  assign n11174 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:40  */
  assign n11175 = csr[11:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:54  */
  assign n11177 = n11175 == 5'b10111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:27  */
  assign n11178 = n11177 & n11174;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1932:21  */
  assign n11179 = csr[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1932:34  */
  assign n11181 = n11179 == 4'b0010;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:84  */
  assign n11182 = n11181 & n11178;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1933:28  */
  assign n11183 = csr[79:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:57  */
  assign n11184 = cnt[143:112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:80  */
  assign n11185 = cnt[307]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:62  */
  assign n11186 = {31'b0, n11185};  //  uext
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1935:62  */
  assign n11187 = n11184 + n11186;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1931:9  */
  assign n11188 = n11182 ? n11183 : n11187;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:58  */
  assign n11199 = cnt[47:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:50  */
  assign n11201 = {1'b0, n11199};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:81  */
  assign n11202 = cnt[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:63  */
  assign n11203 = {32'b0, n11202};  //  uext
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1941:63  */
  assign n11204 = n11201 + n11203;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1952:29  */
  assign n11206 = cnt[111:80]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1953:29  */
  assign n11209 = cnt[207:176]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1954:29  */
  assign n11212 = cnt[47:16]; // extract
  assign n11213 = n11207[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1955:29  */
  assign n11214 = cnt[143:112]; // extract
  assign n11215 = n11210[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2018:16  */
  assign n11220 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2022:42  */
  assign n11223 = cnt_event[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2022:88  */
  assign n11224 = csr[306]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2022:67  */
  assign n11225 = ~n11224;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2022:62  */
  assign n11226 = n11223 & n11225;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2022:113  */
  assign n11227 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2022:98  */
  assign n11228 = ~n11227;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2022:93  */
  assign n11229 = n11226 & n11228;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2024:42  */
  assign n11231 = cnt_event[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2024:88  */
  assign n11232 = csr[308]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2024:67  */
  assign n11233 = ~n11232;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2024:62  */
  assign n11234 = n11231 & n11233;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2024:113  */
  assign n11235 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2024:98  */
  assign n11236 = ~n11235;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2024:93  */
  assign n11237 = n11234 & n11236;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11239 = hpmevent_cfg[155:144]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11240 = cnt_event & n11239;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11246 = n11240[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11248 = 1'b0 | n11246;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11250 = n11240[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11251 = n11248 | n11250;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11252 = n11240[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11253 = n11251 | n11252;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11254 = n11240[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11255 = n11253 | n11254;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11256 = n11240[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11257 = n11255 | n11256;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11258 = n11240[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11259 = n11257 | n11258;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11260 = n11240[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11261 = n11259 | n11260;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11262 = n11240[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11263 = n11261 | n11262;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11264 = n11240[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11265 = n11263 | n11264;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11266 = n11240[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11267 = n11265 | n11266;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11268 = n11240[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11269 = n11267 | n11268;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11270 = n11240[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11271 = n11269 | n11270;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11272 = csr[309]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11273 = ~n11272;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11274 = n11271 & n11273;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11275 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11276 = ~n11275;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11277 = n11274 & n11276;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11279 = hpmevent_cfg[143:132]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11280 = cnt_event & n11279;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11286 = n11280[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11288 = 1'b0 | n11286;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11290 = n11280[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11291 = n11288 | n11290;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11292 = n11280[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11293 = n11291 | n11292;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11294 = n11280[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11295 = n11293 | n11294;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11296 = n11280[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11297 = n11295 | n11296;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11298 = n11280[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11299 = n11297 | n11298;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11300 = n11280[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11301 = n11299 | n11300;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11302 = n11280[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11303 = n11301 | n11302;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11304 = n11280[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11305 = n11303 | n11304;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11306 = n11280[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11307 = n11305 | n11306;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11308 = n11280[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11309 = n11307 | n11308;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11310 = n11280[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11311 = n11309 | n11310;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11312 = csr[310]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11313 = ~n11312;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11314 = n11311 & n11313;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11315 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11316 = ~n11315;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11317 = n11314 & n11316;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11319 = hpmevent_cfg[131:120]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11320 = cnt_event & n11319;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11326 = n11320[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11328 = 1'b0 | n11326;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11330 = n11320[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11331 = n11328 | n11330;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11332 = n11320[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11333 = n11331 | n11332;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11334 = n11320[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11335 = n11333 | n11334;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11336 = n11320[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11337 = n11335 | n11336;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11338 = n11320[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11339 = n11337 | n11338;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11340 = n11320[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11341 = n11339 | n11340;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11342 = n11320[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11343 = n11341 | n11342;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11344 = n11320[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11345 = n11343 | n11344;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11346 = n11320[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11347 = n11345 | n11346;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11348 = n11320[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11349 = n11347 | n11348;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11350 = n11320[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11351 = n11349 | n11350;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11352 = csr[311]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11353 = ~n11352;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11354 = n11351 & n11353;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11355 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11356 = ~n11355;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11357 = n11354 & n11356;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11359 = hpmevent_cfg[119:108]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11360 = cnt_event & n11359;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11366 = n11360[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11368 = 1'b0 | n11366;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11370 = n11360[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11371 = n11368 | n11370;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11372 = n11360[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11373 = n11371 | n11372;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11374 = n11360[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11375 = n11373 | n11374;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11376 = n11360[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11377 = n11375 | n11376;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11378 = n11360[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11379 = n11377 | n11378;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11380 = n11360[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11381 = n11379 | n11380;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11382 = n11360[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11383 = n11381 | n11382;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11384 = n11360[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11385 = n11383 | n11384;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11386 = n11360[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11387 = n11385 | n11386;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11388 = n11360[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11389 = n11387 | n11388;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11390 = n11360[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11391 = n11389 | n11390;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11392 = csr[312]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11393 = ~n11392;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11394 = n11391 & n11393;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11395 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11396 = ~n11395;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11397 = n11394 & n11396;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11399 = hpmevent_cfg[107:96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11400 = cnt_event & n11399;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11406 = n11400[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11408 = 1'b0 | n11406;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11410 = n11400[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11411 = n11408 | n11410;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11412 = n11400[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11413 = n11411 | n11412;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11414 = n11400[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11415 = n11413 | n11414;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11416 = n11400[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11417 = n11415 | n11416;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11418 = n11400[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11419 = n11417 | n11418;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11420 = n11400[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11421 = n11419 | n11420;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11422 = n11400[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11423 = n11421 | n11422;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11424 = n11400[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11425 = n11423 | n11424;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11426 = n11400[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11427 = n11425 | n11426;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11428 = n11400[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11429 = n11427 | n11428;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11430 = n11400[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11431 = n11429 | n11430;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11432 = csr[313]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11433 = ~n11432;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11434 = n11431 & n11433;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11435 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11436 = ~n11435;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11437 = n11434 & n11436;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11439 = hpmevent_cfg[95:84]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11440 = cnt_event & n11439;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11446 = n11440[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11448 = 1'b0 | n11446;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11450 = n11440[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11451 = n11448 | n11450;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11452 = n11440[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11453 = n11451 | n11452;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11454 = n11440[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11455 = n11453 | n11454;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11456 = n11440[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11457 = n11455 | n11456;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11458 = n11440[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11459 = n11457 | n11458;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11460 = n11440[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11461 = n11459 | n11460;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11462 = n11440[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11463 = n11461 | n11462;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11464 = n11440[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11465 = n11463 | n11464;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11466 = n11440[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11467 = n11465 | n11466;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11468 = n11440[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11469 = n11467 | n11468;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11470 = n11440[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11471 = n11469 | n11470;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11472 = csr[314]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11473 = ~n11472;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11474 = n11471 & n11473;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11475 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11476 = ~n11475;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11477 = n11474 & n11476;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11479 = hpmevent_cfg[83:72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11480 = cnt_event & n11479;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11486 = n11480[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11488 = 1'b0 | n11486;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11490 = n11480[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11491 = n11488 | n11490;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11492 = n11480[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11493 = n11491 | n11492;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11494 = n11480[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11495 = n11493 | n11494;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11496 = n11480[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11497 = n11495 | n11496;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11498 = n11480[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11499 = n11497 | n11498;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11500 = n11480[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11501 = n11499 | n11500;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11502 = n11480[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11503 = n11501 | n11502;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11504 = n11480[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11505 = n11503 | n11504;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11506 = n11480[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11507 = n11505 | n11506;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11508 = n11480[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11509 = n11507 | n11508;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11510 = n11480[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11511 = n11509 | n11510;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11512 = csr[315]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11513 = ~n11512;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11514 = n11511 & n11513;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11515 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11516 = ~n11515;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11517 = n11514 & n11516;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11519 = hpmevent_cfg[71:60]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11520 = cnt_event & n11519;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11526 = n11520[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11528 = 1'b0 | n11526;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11530 = n11520[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11531 = n11528 | n11530;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11532 = n11520[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11533 = n11531 | n11532;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11534 = n11520[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11535 = n11533 | n11534;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11536 = n11520[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11537 = n11535 | n11536;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11538 = n11520[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11539 = n11537 | n11538;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11540 = n11520[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11541 = n11539 | n11540;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11542 = n11520[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11543 = n11541 | n11542;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11544 = n11520[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11545 = n11543 | n11544;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11546 = n11520[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11547 = n11545 | n11546;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11548 = n11520[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11549 = n11547 | n11548;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11550 = n11520[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11551 = n11549 | n11550;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11552 = csr[316]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11553 = ~n11552;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11554 = n11551 & n11553;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11555 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11556 = ~n11555;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11557 = n11554 & n11556;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11559 = hpmevent_cfg[59:48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11560 = cnt_event & n11559;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11566 = n11560[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11568 = 1'b0 | n11566;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11570 = n11560[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11571 = n11568 | n11570;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11572 = n11560[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11573 = n11571 | n11572;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11574 = n11560[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11575 = n11573 | n11574;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11576 = n11560[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11577 = n11575 | n11576;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11578 = n11560[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11579 = n11577 | n11578;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11580 = n11560[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11581 = n11579 | n11580;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11582 = n11560[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11583 = n11581 | n11582;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11584 = n11560[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11585 = n11583 | n11584;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11586 = n11560[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11587 = n11585 | n11586;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11588 = n11560[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11589 = n11587 | n11588;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11590 = n11560[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11591 = n11589 | n11590;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11592 = csr[317]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11593 = ~n11592;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11594 = n11591 & n11593;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11595 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11596 = ~n11595;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11597 = n11594 & n11596;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11599 = hpmevent_cfg[47:36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11600 = cnt_event & n11599;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11606 = n11600[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11608 = 1'b0 | n11606;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11610 = n11600[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11611 = n11608 | n11610;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11612 = n11600[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11613 = n11611 | n11612;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11614 = n11600[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11615 = n11613 | n11614;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11616 = n11600[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11617 = n11615 | n11616;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11618 = n11600[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11619 = n11617 | n11618;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11620 = n11600[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11621 = n11619 | n11620;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11622 = n11600[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11623 = n11621 | n11622;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11624 = n11600[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11625 = n11623 | n11624;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11626 = n11600[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11627 = n11625 | n11626;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11628 = n11600[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11629 = n11627 | n11628;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11630 = n11600[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11631 = n11629 | n11630;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11632 = csr[318]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11633 = ~n11632;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11634 = n11631 & n11633;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11635 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11636 = ~n11635;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11637 = n11634 & n11636;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11639 = hpmevent_cfg[35:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11640 = cnt_event & n11639;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11646 = n11640[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11648 = 1'b0 | n11646;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11650 = n11640[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11651 = n11648 | n11650;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11652 = n11640[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11653 = n11651 | n11652;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11654 = n11640[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11655 = n11653 | n11654;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11656 = n11640[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11657 = n11655 | n11656;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11658 = n11640[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11659 = n11657 | n11658;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11660 = n11640[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11661 = n11659 | n11660;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11662 = n11640[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11663 = n11661 | n11662;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11664 = n11640[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11665 = n11663 | n11664;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11666 = n11640[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11667 = n11665 | n11666;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11668 = n11640[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11669 = n11667 | n11668;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11670 = n11640[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11671 = n11669 | n11670;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11672 = csr[319]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11673 = ~n11672;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11674 = n11671 & n11673;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11675 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11676 = ~n11675;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11677 = n11674 & n11676;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11679 = hpmevent_cfg[23:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11680 = cnt_event & n11679;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11686 = n11680[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11688 = 1'b0 | n11686;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11690 = n11680[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11691 = n11688 | n11690;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11692 = n11680[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11693 = n11691 | n11692;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11694 = n11680[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11695 = n11693 | n11694;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11696 = n11680[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11697 = n11695 | n11696;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11698 = n11680[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11699 = n11697 | n11698;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11700 = n11680[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11701 = n11699 | n11700;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11702 = n11680[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11703 = n11701 | n11702;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11704 = n11680[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11705 = n11703 | n11704;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11706 = n11680[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11707 = n11705 | n11706;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11708 = n11680[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11709 = n11707 | n11708;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11710 = n11680[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11711 = n11709 | n11710;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11712 = csr[320]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11713 = ~n11712;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11714 = n11711 & n11713;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11715 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11716 = ~n11715;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11717 = n11714 & n11716;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:73  */
  assign n11719 = hpmevent_cfg[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:57  */
  assign n11720 = cnt_event & n11719;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11726 = n11720[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11728 = 1'b0 | n11726;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11730 = n11720[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11731 = n11728 | n11730;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11732 = n11720[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11733 = n11731 | n11732;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11734 = n11720[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11735 = n11733 | n11734;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11736 = n11720[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11737 = n11735 | n11736;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11738 = n11720[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11739 = n11737 | n11738;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11740 = n11720[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11741 = n11739 | n11740;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11742 = n11720[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11743 = n11741 | n11742;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11744 = n11720[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11745 = n11743 | n11744;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11746 = n11720[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11747 = n11745 | n11746;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11748 = n11720[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11749 = n11747 | n11748;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n11750 = n11720[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n11751 = n11749 | n11750;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:104  */
  assign n11752 = csr[321]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:83  */
  assign n11753 = ~n11752;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:78  */
  assign n11754 = n11751 & n11753;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:129  */
  assign n11755 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:114  */
  assign n11756 = ~n11755;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2027:109  */
  assign n11757 = n11754 & n11756;
  assign n11758 = {n11757, n11717, n11677, n11637, n11597, n11557, n11517, n11477, n11437, n11397, n11357, n11317, n11277, n11237, 1'b0, n11229};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2033:56  */
  assign n11764 = ~sleep_mode;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2033:39  */
  assign n11765 = n11764 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2035:56  */
  assign n11769 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2035:62  */
  assign n11771 = n11769 == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2035:39  */
  assign n11772 = n11771 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2038:62  */
  assign n11775 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2038:68  */
  assign n11777 = n11775 == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2038:99  */
  assign n11778 = exe_engine[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2038:83  */
  assign n11779 = n11778 & n11777;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2038:45  */
  assign n11780 = n11779 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2039:62  */
  assign n11783 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2039:68  */
  assign n11785 = n11783 == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2039:101  */
  assign n11786 = issue_engine[86:85]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2039:107  */
  assign n11788 = n11786 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2039:83  */
  assign n11789 = n11788 & n11785;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2039:45  */
  assign n11790 = n11789 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2040:62  */
  assign n11793 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2040:68  */
  assign n11795 = n11793 == 4'b0110;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2040:45  */
  assign n11796 = n11795 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2041:62  */
  assign n11799 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2041:68  */
  assign n11801 = n11799 == 4'b0111;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2041:45  */
  assign n11802 = n11801 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2042:62  */
  assign n11805 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2042:68  */
  assign n11807 = n11805 == 4'b1000;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2042:45  */
  assign n11808 = n11807 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2043:56  */
  assign n11811 = ctrl[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2043:83  */
  assign n11812 = opcode[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2043:87  */
  assign n11813 = ~n11812;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2043:104  */
  assign n11814 = opcode[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2043:94  */
  assign n11815 = n11813 | n11814;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2043:71  */
  assign n11816 = n11815 & n11811;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2043:45  */
  assign n11817 = n11816 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2044:56  */
  assign n11820 = ctrl[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2044:83  */
  assign n11821 = opcode[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2044:104  */
  assign n11822 = opcode[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2044:94  */
  assign n11823 = n11821 | n11822;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2044:71  */
  assign n11824 = n11823 & n11820;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2044:45  */
  assign n11825 = n11824 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2045:56  */
  assign n11828 = ctrl[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2045:64  */
  assign n11829 = ~n11828;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2045:87  */
  assign n11830 = exe_engine[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2045:93  */
  assign n11832 = n11830 == 4'b1011;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2045:71  */
  assign n11833 = n11832 & n11829;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2045:45  */
  assign n11834 = n11833 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2046:61  */
  assign n11837 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2046:45  */
  assign n11838 = n11837 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2060:18  */
  assign n11841 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2063:24  */
  assign n11844 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2063:28  */
  assign n11845 = ~n11844;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2064:25  */
  assign n11846 = trap_ctrl[97]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2064:62  */
  assign n11847 = trap_ctrl[62]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2064:42  */
  assign n11848 = n11847 & n11846;
  assign n11850 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2064:11  */
  assign n11851 = n11848 ? 1'b1 : n11850;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2068:25  */
  assign n11852 = trap_ctrl[99]; // extract
  assign n11854 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2068:11  */
  assign n11855 = n11852 ? 1'b0 : n11854;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2063:9  */
  assign n11856 = n11845 ? n11851 : n11855;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2076:40  */
  assign n11861 = trap_ctrl[106]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2076:67  */
  assign n11862 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2076:52  */
  assign n11863 = ~n11862;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2076:47  */
  assign n11864 = n11861 & n11863;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2076:80  */
  assign n11865 = csr[426]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2076:72  */
  assign n11866 = n11864 & n11865;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2076:102  */
  assign n11867 = csr[427]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2076:94  */
  assign n11868 = n11866 & n11867;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2077:40  */
  assign n11869 = trap_ctrl[105]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2077:63  */
  assign n11870 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2078:40  */
  assign n11871 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2078:59  */
  assign n11872 = csr[322]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2078:51  */
  assign n11873 = n11871 & n11872;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2077:67  */
  assign n11874 = n11870 | n11873;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2079:40  */
  assign n11875 = csr[136]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2079:32  */
  assign n11876 = ~n11875;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2079:59  */
  assign n11877 = csr[323]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2079:51  */
  assign n11878 = n11876 & n11877;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2078:73  */
  assign n11879 = n11874 | n11878;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2077:47  */
  assign n11880 = n11869 & n11879;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2080:64  */
  assign n11881 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2080:49  */
  assign n11882 = ~n11881;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2080:44  */
  assign n11883 = irq_dbg_i & n11882;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2081:34  */
  assign n11884 = csr[324]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2081:64  */
  assign n11885 = debug_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2081:49  */
  assign n11886 = ~n11885;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2081:44  */
  assign n11887 = n11884 & n11886;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2100:36  */
  assign n11890 = csr[322]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2103:36  */
  assign n11893 = csr[323]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2103:49  */
  assign n11895 = 1'b1 ? n11893 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2107:36  */
  assign n11900 = csr[328:326]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2111:36  */
  assign n11904 = csr[324]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2112:47  */
  assign n11905 = csr[325]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2112:47  */
  assign n11906 = csr[325]; // extract
  assign n11907 = {n11905, n11906};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2122:39  */
  assign n11909 = csr[425]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2123:52  */
  assign n11910 = ~hw_trigger_fired;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2122:61  */
  assign n11911 = n11910 & n11909;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2124:45  */
  assign n11912 = csr[491:461]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2124:79  */
  assign n11913 = exe_engine[100:70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2124:63  */
  assign n11914 = n11912 == n11913;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2123:59  */
  assign n11915 = n11914 & n11911;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2122:29  */
  assign n11916 = n11915 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2130:18  */
  assign n11919 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2133:30  */
  assign n11921 = ~hw_trigger_fired;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2134:69  */
  assign n11922 = trap_ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2134:48  */
  assign n11923 = hw_trigger_match & n11922;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2135:20  */
  assign n11924 = csr[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2135:39  */
  assign n11925 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2135:44  */
  assign n11927 = n11925 == 12'b011110100001;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2135:30  */
  assign n11928 = n11927 & n11924;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2135:74  */
  assign n11929 = csr[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2135:79  */
  assign n11930 = ~n11929;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2135:60  */
  assign n11931 = n11930 & n11928;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2135:9  */
  assign n11933 = n11931 ? 1'b0 : hw_trigger_fired;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2133:9  */
  assign n11934 = n11921 ? n11923 : n11933;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2154:38  */
  assign n11940 = csr[427]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2163:46  */
  assign n11948 = csr[426]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2163:40  */
  assign n11950 = {3'b000, n11948};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2170:38  */
  assign n11958 = csr[425]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:313:5  */
  always @(posedge clk_i or posedge n7435)
    if (n7435)
      n11961 <= 1'b0;
    else
      n11961 <= n7493;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:313:5  */
  always @(posedge clk_i or posedge n7435)
    if (n7435)
      n11962 <= n7499;
    else
      n11962 <= n7494;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:308:5  */
  assign n11963 = {n11961, n7518, n8307, n11962};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:308:5  */
  assign n11964 = {\prefetch_buffer_n2_prefetch_buffer_inst.avail_o , \prefetch_buffer_n1_prefetch_buffer_inst.avail_o , \prefetch_buffer_n2_prefetch_buffer_inst.free_o , \prefetch_buffer_n1_prefetch_buffer_inst.free_o , n7678, n7675, n7544, n7536, \prefetch_buffer_n1_prefetch_buffer_inst.rdata_o , \prefetch_buffer_n2_prefetch_buffer_inst.rdata_o , n7521, n7524};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:423:7  */
  always @(posedge clk_i or posedge n7570)
    if (n7570)
      n11965 <= 1'b0;
    else
      n11965 <= n7584;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:421:7  */
  assign n11966 = {n8308, n7664, \issue_engine_enabled_neorv32_cpu_decompressor_inst.instr_o , n7671, n7663, n7621, n11965};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:559:5  */
  always @(posedge clk_i or posedge n7817)
    if (n7817)
      n11967 <= n7827;
    else
      n11967 <= exe_engine_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:551:5  */
  assign n11968 = {n8313, n8312, n8311, n8309};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:899:5  */
  always @(posedge clk_i or posedge n8392)
    if (n8392)
      n11969 <= 10'b0000000000;
    else
      n11969 <= n8400;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1298:5  */
  always @(posedge clk_aux_i or posedge n9514)
    if (n9514)
      n11970 <= 1'b0;
    else
      n11970 <= n9528;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1250:5  */
  always @(posedge clk_i or posedge n9341)
    if (n9341)
      n11971 <= 1'b0;
    else
      n11971 <= n9380;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1250:5  */
  always @(posedge clk_i or posedge n9341)
    if (n9341)
      n11972 <= 1'b0;
    else
      n11972 <= n9371;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1197:5  */
  always @(posedge clk_i or posedge n9222)
    if (n9222)
      n11973 <= 7'b0000000;
    else
      n11973 <= n9331;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1149:5  */
  always @(posedge clk_aux_i or posedge n9063)
    if (n9063)
      n11974 <= n9218;
    else
      n11974 <= n9215;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1102:5  */
  always @(posedge clk_i or posedge n8964)
    if (n8964)
      n11975 <= 11'b00000000000;
    else
      n11975 <= n9057;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1100:5  */
  assign n11976 = {n8320, n8319, n8961, n8317, n8316, n9587, n8315, n11971, n8314, n11972, n9338, n11973, n9511, n9497, n9485, n11974, n9420, n11975};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:559:5  */
  always @(posedge clk_i or posedge n7817)
    if (n7817)
      n11977 <= 59'b00000000000000000000000000000000000000000000000000000000000;
    else
      n11977 <= ctrl_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:551:5  */
  assign n11978 = {n8351, n8342, n8352, n7915, n8340, n8338, n8336, n8334, n7869, n8332, n8331, n8330, n8328, n8326, n8346, n8324, n8322};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1650:5  */
  always @(posedge clk_i or posedge n9990)
    if (n9990)
      n11979 <= 32'b00000000000000000000000000000000;
    else
      n11979 <= n11046;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1650:5  */
  always @(posedge clk_i or posedge n9990)
    if (n9990)
      n11980 <= 1'b0;
    else
      n11980 <= n9997;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1386:5  */
  assign n11981 = csr[491:460]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1386:5  */
  assign n11982 = n9960 ? n9805 : n11981;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1386:5  */
  always @(posedge clk_i or posedge n9627)
    if (n9627)
      n11983 <= 32'b00000000000000000000000000000000;
    else
      n11983 <= n11982;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1386:5  */
  always @(posedge clk_i or posedge n9627)
    if (n9627)
      n11984 <= n9978;
    else
      n11984 <= n9965;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1386:5  */
  always @(posedge clk_i or posedge n9627)
    if (n9627)
      n11985 <= n9977;
    else
      n11985 <= n9964;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1386:5  */
  always @(posedge clk_i or posedge n9627)
    if (n9627)
      n11986 <= n9976;
    else
      n11986 <= n9963;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1386:5  */
  always @(posedge clk_i or posedge n9627)
    if (n9627)
      n11987 <= 1'b0;
    else
      n11987 <= n9663;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1323:5  */
  assign n11988 = csr[11:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1323:5  */
  assign n11989 = n9593 ? n9594 : n11988;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1323:5  */
  always @(posedge clk_i or posedge n9589)
    if (n9589)
      n11990 <= 12'b000000000000;
    else
      n11990 <= n11989;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1321:5  */
  assign n11991 = {n11983, 4'b0110, n11940, 1'b0, 1'b0, 1'b0, 1'b0, hw_trigger_fired, 1'b0, 2'b00, 3'b000, n11950, 1'b0, 4'b0000, 1'b1, 1'b0, 1'b0, 1'b1, n11958, 1'b0, 1'b0, n11984, 4'b0100, 12'b000000000000, n11890, 1'b0, 1'b0, n11895, 1'b0, 1'b1, 1'b0, n11900, 1'b0, 1'b1, 1'b0, n11904, n11907, n11985, n9987, n11986, n11979, n9621, n9603, n8354, n11980, n8353, n11987, n11990};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2020:5  */
  always @(posedge clk_i or posedge n11220)
    if (n11220)
      n11992 <= 16'b0000000000000000;
    else
      n11992 <= n11758;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11156)
    if (n11156)
      n11993 <= 1'b0;
    else
      n11993 <= n11173;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11156)
    if (n11156)
      n11994 <= 32'b00000000000000000000000000000000;
    else
      n11994 <= n11188;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11156)
    if (n11156)
      n11995 <= 32'b00000000000000000000000000000000;
    else
      n11995 <= n11172;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11106)
    if (n11106)
      n11996 <= 1'b0;
    else
      n11996 <= n11123;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11106)
    if (n11106)
      n11997 <= 32'b00000000000000000000000000000000;
    else
      n11997 <= n11138;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11106)
    if (n11106)
      n11998 <= 32'b00000000000000000000000000000000;
    else
      n11998 <= n11122;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11056)
    if (n11056)
      n11999 <= 1'b0;
    else
      n11999 <= n11073;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11056)
    if (n11056)
      n12000 <= 32'b00000000000000000000000000000000;
    else
      n12000 <= n11088;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1919:7  */
  always @(posedge clk_i or posedge n11056)
    if (n11056)
      n12001 <= 32'b00000000000000000000000000000000;
    else
      n12001 <= n11072;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:7  */
  assign n12002 = {n11999, n11996, n11993, n11104, n11154, n11204, n12000, n11997, n11994, n12001, n11998, n11995, n11992};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:7  */
  assign n12003 = {n11209, n11215, n11214};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:7  */
  assign n12004 = {n11206, n11213, n11212};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:7  */
  assign n12005 = {n11838, n11834, n11825, n11817, n11808, n11802, n11796, n11790, n11780, n11772, 1'b0, n11765};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2062:7  */
  always @(posedge clk_i or posedge n11841)
    if (n11841)
      n12006 <= 1'b0;
    else
      n12006 <= n11856;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2060:7  */
  assign n12007 = {n11887, n11883, n11880, n11868, n12006};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:7  */
  assign n12008 = {n8731, n8749, n8792};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2132:7  */
  always @(posedge clk_i or posedge n11919)
    if (n11919)
      n12009 <= 1'b0;
    else
      n12009 <= n11934;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:2130:7  */
  assign n12010 = {n8390, n8389, sleep_mode, n8388, opcode, n8387, n8386, n8384, n8381, n8379, n8374, n8373, n8372, n8371, n8370, n8369, n8368, n8367, n8366, n8365, n8364, n8363, n8362, n8361, n8360, n8356};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:1915:7  */
  assign n12011 = {n7554, sleep_mode, n7553, 4'b0000, 1'b0, n7546, 1'b1, 1'b0, n7514, 4'b0000, 32'b00000000000000000000000000000000, n7505};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu_control.vhd:503:5  */
  always @(posedge clk_i or posedge n7680)
    if (n7680)
      n12012 <= 32'b00000000000000000000000000000000;
    else
      n12012 <= n7796;
endmodule

module neorv32_debug_dm_1_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk_i,
   input  rstn_i,
   input  [6:0] \dmi_req_i_dmi_req_i[addr] ,
   input  [1:0] \dmi_req_i_dmi_req_i[op] ,
   input  [31:0] \dmi_req_i_dmi_req_i[data] ,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   output [31:0] \dmi_rsp_o_dmi_rsp_o[data] ,
   output \dmi_rsp_o_dmi_rsp_o[ack] ,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output ndmrstn_o,
   output halt_req_o);
  wire [40:0] n6239;
  wire [31:0] n6241;
  wire n6242;
  wire [79:0] n6243;
  wire [31:0] n6245;
  wire n6246;
  wire n6247;
  wire dmi_wren;
  wire dmi_wren_auth;
  wire dmi_rden;
  wire dmi_rden_auth;
  wire [113:0] dm_reg;
  wire [127:0] cpu_progbuf;
  wire [45:0] dm_ctrl;
  wire [35:0] auth;
  wire accen;
  wire rden;
  wire wren;
  wire cpu_rsp_dec;
  wire [38:0] dci;
  wire [1:0] n6251;
  wire n6253;
  wire n6254;
  wire [1:0] n6257;
  wire n6259;
  wire n6260;
  wire n6263;
  wire n6266;
  wire n6269;
  wire n6278;
  wire n6279;
  localparam [31:0] n6281 = 32'b00000000000000000010000000100011;
  wire [2:0] n6290;
  wire [6:0] n6291;
  wire n6293;
  wire [2:0] n6294;
  wire n6296;
  wire [2:0] n6298;
  wire [2:0] n6299;
  wire n6301;
  wire n6302;
  wire n6303;
  wire n6304;
  wire [2:0] n6306;
  wire [2:0] n6307;
  wire [2:0] n6308;
  wire n6310;
  wire [7:0] n6311;
  wire n6313;
  wire n6314;
  wire n6315;
  wire n6316;
  wire [2:0] n6317;
  wire n6319;
  wire n6320;
  wire n6321;
  wire n6322;
  wire n6323;
  wire n6324;
  wire n6325;
  wire [10:0] n6326;
  wire n6328;
  wire n6329;
  wire n6330;
  wire n6332;
  wire n6333;
  wire n6334;
  wire n6341;
  wire [2:0] n6346;
  wire n6347;
  wire [2:0] n6350;
  wire n6351;
  wire n6352;
  wire n6354;
  wire n6355;
  wire n6356;
  wire n6357;
  wire [4:0] n6360;
  wire [7:0] n6363;
  wire [6:0] n6364;
  localparam [31:0] n6365 = 32'b00000000000000000010000000000011;
  wire [4:0] n6368;
  wire [7:0] n6369;
  wire [6:0] n6370;
  wire [31:0] n6371;
  wire [31:0] n6372;
  wire [31:0] n6373;
  wire [31:0] n6375;
  wire n6376;
  wire n6379;
  wire n6380;
  wire n6382;
  wire n6383;
  wire n6384;
  wire n6391;
  wire [2:0] n6394;
  wire [2:0] n6395;
  wire n6397;
  wire n6399;
  wire n6400;
  wire n6401;
  wire n6408;
  wire [2:0] n6411;
  wire [2:0] n6412;
  wire n6414;
  wire n6417;
  wire [5:0] n6419;
  reg [2:0] n6420;
  wire [31:0] n6421;
  reg [31:0] n6422;
  wire n6423;
  reg n6424;
  reg n6425;
  reg n6426;
  reg n6427;
  wire [2:0] n6428;
  wire n6430;
  wire n6431;
  wire n6433;
  wire n6435;
  wire n6437;
  wire n6438;
  wire n6439;
  wire [2:0] n6441;
  wire [2:0] n6442;
  wire [2:0] n6443;
  wire [2:0] n6444;
  wire [2:0] n6445;
  wire n6446;
  wire [2:0] n6448;
  wire [2:0] n6449;
  wire [2:0] n6450;
  wire [37:0] n6451;
  wire [37:0] n6452;
  wire [2:0] n6453;
  wire [37:0] n6454;
  wire n6455;
  wire [37:0] n6462;
  wire [2:0] n6468;
  wire n6470;
  wire n6471;
  wire n6474;
  wire n6480;
  wire n6482;
  wire n6484;
  wire n6486;
  wire n6487;
  wire n6488;
  wire n6489;
  wire n6490;
  wire n6492;
  wire n6493;
  wire n6494;
  wire n6496;
  wire n6498;
  wire n6499;
  wire n6500;
  wire n6501;
  wire n6502;
  wire n6504;
  wire n6506;
  wire n6507;
  wire n6508;
  wire n6510;
  wire n6511;
  wire n6512;
  wire n6513;
  wire n6514;
  wire n6516;
  wire n6517;
  wire n6518;
  wire n6520;
  wire n6521;
  wire n6522;
  wire [3:0] n6523;
  wire [3:0] n6526;
  wire n6530;
  wire [6:0] n6550;
  wire n6552;
  wire n6553;
  wire n6554;
  wire n6555;
  wire [2:0] n6556;
  wire n6557;
  wire [5:0] n6558;
  wire n6559;
  wire n6560;
  wire n6561;
  wire [2:0] n6562;
  wire [5:0] n6563;
  wire [5:0] n6564;
  wire n6565;
  wire n6566;
  wire n6567;
  wire [1:0] n6568;
  wire [1:0] n6569;
  wire [1:0] n6570;
  wire n6571;
  wire [2:0] n6572;
  wire [5:0] n6573;
  wire [5:0] n6574;
  wire [6:0] n6575;
  wire n6577;
  wire n6578;
  wire n6579;
  wire n6580;
  wire n6581;
  wire [2:0] n6582;
  wire n6584;
  wire n6585;
  wire [31:0] n6586;
  wire [31:0] n6587;
  wire [31:0] n6588;
  wire [6:0] n6589;
  wire n6591;
  wire n6592;
  wire n6593;
  wire n6594;
  wire n6595;
  wire n6596;
  wire n6597;
  wire n6598;
  wire [2:0] n6599;
  wire [2:0] n6600;
  wire [2:0] n6601;
  wire [6:0] n6602;
  wire n6604;
  wire n6605;
  wire n6606;
  wire [6:0] n6607;
  wire n6609;
  wire n6610;
  wire n6611;
  wire n6612;
  wire [6:0] n6613;
  wire n6615;
  wire n6616;
  wire n6617;
  wire n6618;
  wire n6620;
  wire n6621;
  wire [6:0] n6622;
  wire n6624;
  wire n6625;
  wire [2:0] n6626;
  wire n6628;
  wire n6629;
  wire n6631;
  wire [6:0] n6632;
  wire n6634;
  wire n6635;
  wire n6636;
  wire n6637;
  wire n6638;
  wire [31:0] n6639;
  wire [31:0] n6640;
  wire [31:0] n6641;
  wire [6:0] n6642;
  wire n6644;
  wire n6645;
  wire n6646;
  wire n6647;
  wire n6648;
  wire [31:0] n6649;
  wire [31:0] n6650;
  wire [31:0] n6651;
  wire n6652;
  wire n6653;
  wire [6:0] n6654;
  wire n6656;
  wire [6:0] n6657;
  wire n6659;
  wire n6660;
  wire [6:0] n6661;
  wire n6663;
  wire n6664;
  wire [6:0] n6665;
  wire n6667;
  wire n6668;
  wire [6:0] n6669;
  wire n6671;
  wire n6672;
  wire [6:0] n6673;
  wire n6675;
  wire n6676;
  wire n6677;
  wire n6679;
  wire [106:0] n6680;
  wire [1:0] n6681;
  wire [106:0] n6688;
  wire [1:0] n6689;
  wire n6695;
  wire n6696;
  wire [1:0] n6697;
  wire n6699;
  wire n6700;
  wire n6701;
  wire [2:0] n6704;
  wire n6706;
  wire n6707;
  wire [6:0] n6710;
  wire n6712;
  wire n6713;
  wire n6714;
  wire n6715;
  wire n6716;
  wire n6717;
  wire n6719;
  wire n6720;
  wire n6721;
  wire n6722;
  wire n6723;
  wire n6725;
  wire n6727;
  wire n6729;
  wire n6730;
  wire n6731;
  wire n6733;
  wire n6734;
  wire [31:0] n6736;
  wire n6737;
  wire n6738;
  wire [31:0] n6739;
  wire [31:0] n6740;
  wire n6741;
  wire n6742;
  wire [31:0] n6743;
  wire [31:0] n6744;
  wire n6747;
  wire n6753;
  localparam [31:0] n6754 = 32'b00000000000000000000000000000000;
  wire [6:0] n6755;
  localparam [8:0] n6756 = 9'b000000000;
  wire n6760;
  wire n6761;
  wire n6762;
  wire n6769;
  wire n6772;
  wire n6773;
  wire n6774;
  wire n6781;
  wire n6784;
  wire n6785;
  wire n6786;
  wire n6793;
  wire n6796;
  wire n6797;
  wire n6798;
  wire n6805;
  wire n6807;
  wire n6808;
  wire n6809;
  wire n6810;
  wire n6812;
  wire n6813;
  wire n6814;
  wire n6821;
  wire n6823;
  wire n6825;
  wire n6826;
  wire n6827;
  wire n6834;
  wire n6836;
  wire n6838;
  wire n6839;
  wire n6840;
  wire n6847;
  wire n6850;
  wire n6851;
  wire n6852;
  wire n6859;
  wire n6863;
  wire n6864;
  localparam [3:0] n6865 = 4'b0011;
  wire n6867;
  wire [2:0] n6874;
  wire [9:0] n6876;
  localparam [9:0] n6877 = 10'b0000000000;
  localparam [1:0] n6878 = 2'b00;
  wire n6881;
  wire n6882;
  wire n6884;
  localparam [7:0] n6885 = 8'b00000000;
  localparam [3:0] n6886 = 4'b0001;
  localparam [2:0] n6887 = 3'b000;
  localparam [3:0] n6889 = 4'b0001;
  localparam [11:0] n6890 = 12'b111100000000;
  wire n6892;
  localparam [7:0] n6893 = 8'b00000000;
  localparam [4:0] n6894 = 5'b00010;
  wire [2:0] n6895;
  wire n6896;
  wire [2:0] n6898;
  localparam [3:0] n6899 = 4'b0000;
  localparam [3:0] n6900 = 4'b0001;
  wire n6902;
  wire n6903;
  wire n6904;
  wire n6905;
  wire n6907;
  wire [31:0] n6908;
  wire n6910;
  wire [31:0] n6911;
  wire n6913;
  wire n6914;
  wire n6916;
  localparam [31:0] n6917 = 32'b00000000000000000000000000000000;
  wire [7:0] n6918;
  wire n6919;
  wire n6920;
  wire n6921;
  wire n6922;
  wire n6923;
  wire n6924;
  reg n6925;
  wire n6926;
  wire n6927;
  wire n6928;
  wire n6929;
  wire n6930;
  wire n6931;
  wire n6932;
  reg n6933;
  wire n6934;
  wire n6935;
  wire n6936;
  wire n6937;
  wire n6938;
  wire n6939;
  wire n6940;
  reg n6941;
  wire n6942;
  wire n6943;
  wire n6944;
  wire n6945;
  wire n6946;
  wire n6947;
  wire n6948;
  reg n6949;
  wire n6950;
  wire n6951;
  wire n6952;
  wire n6953;
  wire n6954;
  wire n6955;
  wire n6956;
  reg n6957;
  wire n6958;
  wire n6959;
  wire n6960;
  wire n6961;
  wire n6962;
  wire n6963;
  wire n6964;
  reg n6965;
  wire n6966;
  wire n6967;
  wire n6968;
  wire n6969;
  wire n6970;
  wire n6971;
  wire n6972;
  reg n6973;
  wire n6974;
  wire n6975;
  wire n6976;
  wire n6977;
  wire n6978;
  wire n6979;
  wire n6980;
  reg n6981;
  wire n6982;
  wire n6983;
  wire n6984;
  wire n6985;
  wire n6986;
  wire n6987;
  wire n6988;
  reg n6989;
  wire n6990;
  wire n6991;
  wire n6992;
  wire n6993;
  wire n6994;
  wire n6995;
  wire n6996;
  reg n6997;
  wire n6998;
  wire n6999;
  wire n7000;
  wire n7001;
  wire n7002;
  wire n7003;
  wire n7004;
  reg n7005;
  wire n7006;
  wire n7007;
  wire n7008;
  wire n7009;
  wire n7010;
  wire n7011;
  reg n7012;
  wire n7013;
  wire n7014;
  wire n7015;
  wire n7016;
  wire n7017;
  wire n7018;
  reg n7019;
  wire n7020;
  wire n7021;
  wire n7022;
  wire n7023;
  wire n7024;
  wire n7025;
  reg n7026;
  wire n7027;
  wire n7028;
  wire n7029;
  wire n7030;
  wire n7031;
  wire n7032;
  reg n7033;
  wire n7034;
  wire n7035;
  wire n7036;
  wire n7037;
  wire n7038;
  wire n7039;
  reg n7040;
  wire n7041;
  wire n7042;
  wire n7043;
  wire n7044;
  wire n7045;
  reg n7046;
  wire n7047;
  wire n7048;
  wire n7049;
  wire n7050;
  wire n7051;
  wire n7052;
  reg n7053;
  wire n7054;
  wire n7055;
  wire n7056;
  wire n7057;
  wire n7058;
  wire n7059;
  reg n7060;
  wire n7061;
  wire n7062;
  wire n7063;
  wire n7064;
  wire n7065;
  wire n7066;
  reg n7067;
  wire [1:0] n7068;
  wire [1:0] n7069;
  wire [1:0] n7070;
  wire [1:0] n7071;
  wire [1:0] n7072;
  wire [1:0] n7073;
  reg [1:0] n7074;
  wire n7075;
  wire n7076;
  wire n7077;
  wire n7078;
  wire n7079;
  wire n7080;
  reg n7081;
  wire n7082;
  wire n7083;
  wire n7084;
  wire n7085;
  wire n7086;
  wire n7087;
  wire n7088;
  reg n7089;
  wire [1:0] n7090;
  wire [1:0] n7091;
  wire [1:0] n7092;
  wire [1:0] n7093;
  wire [1:0] n7094;
  wire [1:0] n7095;
  wire [1:0] n7096;
  wire [1:0] n7097;
  reg [1:0] n7098;
  wire n7099;
  wire n7100;
  wire n7101;
  wire n7102;
  wire n7103;
  wire n7104;
  wire n7105;
  reg n7106;
  wire n7107;
  wire n7108;
  wire n7109;
  wire n7110;
  wire n7111;
  wire n7112;
  wire n7113;
  reg n7114;
  wire n7115;
  wire n7116;
  wire n7117;
  wire n7118;
  wire n7119;
  wire n7120;
  wire n7121;
  reg n7122;
  wire n7123;
  wire n7124;
  wire n7125;
  wire n7126;
  wire n7127;
  wire n7128;
  wire n7129;
  reg n7130;
  wire n7131;
  wire n7132;
  wire n7133;
  wire n7134;
  wire n7135;
  wire n7136;
  wire n7137;
  reg n7138;
  wire n7139;
  wire n7140;
  wire n7141;
  wire n7142;
  wire n7143;
  wire n7144;
  wire n7145;
  reg n7146;
  wire n7176;
  wire n7177;
  wire [6:0] n7178;
  wire n7180;
  wire [6:0] n7181;
  wire n7183;
  wire n7184;
  wire [6:0] n7185;
  wire n7187;
  wire n7188;
  wire n7189;
  wire n7192;
  wire [6:0] n7193;
  wire n7195;
  wire n7196;
  wire n7197;
  wire [6:0] n7198;
  wire n7200;
  wire n7201;
  wire n7202;
  wire n7203;
  wire [6:0] n7204;
  wire n7206;
  wire n7207;
  wire n7208;
  wire n7209;
  wire n7210;
  wire n7213;
  wire [32:0] n7214;
  wire [32:0] n7220;
  wire n7226;
  wire n7234;
  wire [31:0] n7235;
  wire [1:0] n7236;
  wire n7238;
  wire n7239;
  wire [31:0] n7240;
  wire [31:0] n7241;
  wire [31:0] n7242;
  wire [31:0] n7243;
  wire [1:0] n7248;
  wire n7250;
  wire n7251;
  wire [1:0] n7252;
  wire n7254;
  wire n7256;
  wire n7258;
  wire [2:0] n7260;
  reg n7261;
  reg n7262;
  reg n7263;
  reg n7264;
  wire [1:0] n7265;
  wire n7266;
  wire n7267;
  wire [1:0] n7268;
  wire [1:0] n7269;
  localparam [31:0] n7270 = 32'b00000000000000000000000000000000;
  wire [1:0] n7271;
  wire [4:0] n7272;
  wire n7280;
  wire [1:0] n7281;
  wire [1:0] n7284;
  wire n7288;
  wire [31:0] n7289;
  wire n7291;
  wire n7292;
  wire n7293;
  wire [2:0] n7294;
  wire n7295;
  wire n7296;
  wire n7297;
  reg n7298;
  wire n7299;
  wire n7300;
  wire n7301;
  reg n7302;
  wire [29:0] n7303;
  wire [29:0] n7304;
  wire [29:0] n7305;
  wire [29:0] n7306;
  reg [29:0] n7307;
  wire [31:0] n7308;
  wire [31:0] n7309;
  wire [33:0] n7310;
  wire [1:0] n7322;
  wire n7328;
  wire n7329;
  wire n7330;
  wire n7331;
  wire n7332;
  wire n7333;
  wire n7334;
  wire n7335;
  wire n7343;
  wire n7345;
  wire n7347;
  wire n7348;
  wire n7349;
  wire n7350;
  wire n7351;
  wire n7352;
  wire n7353;
  reg n7360;
  reg n7361;
  reg [1:0] n7362;
  reg n7363;
  reg [106:0] n7364;
  wire [113:0] n7365;
  wire [127:0] n7366;
  reg [3:0] n7367;
  reg [37:0] n7368;
  reg [2:0] n7369;
  wire [45:0] n7370;
  wire [35:0] n7371;
  reg [31:0] n7372;
  reg [1:0] n7373;
  reg n7374;
  reg n7375;
  reg n7376;
  wire [38:0] n7377;
  reg [32:0] n7378;
  reg [33:0] n7379;
  wire [31:0] n7382; // mem_rd
  wire [31:0] n7383;
  assign \dmi_rsp_o_dmi_rsp_o[data]  = n6241; //(module output)
  assign \dmi_rsp_o_dmi_rsp_o[ack]  = n6242; //(module output)
  assign \bus_rsp_o_bus_rsp_o[data]  = n6245; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n6246; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n6247; //(module output)
  assign ndmrstn_o = n6734; //(module output)
  assign halt_req_o = n6725; //(module output)
  assign n6239 = {\dmi_req_i_dmi_req_i[data] , \dmi_req_i_dmi_req_i[op] , \dmi_req_i_dmi_req_i[addr] };
  assign n6241 = n7378[31:0]; // extract
  assign n6242 = n7378[32]; // extract
  assign n6243 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:256:3  */
  assign n6245 = n7379[31:0]; // extract
  assign n6246 = n7379[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1152:14  */
  assign n6247 = n7379[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:76:10  */
  assign dmi_wren = n6254; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:76:20  */
  assign dmi_wren_auth = n6263; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:76:35  */
  assign dmi_rden = n6260; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:76:45  */
  assign dmi_rden_auth = n6266; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:100:10  */
  assign dm_reg = n7365; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:104:10  */
  assign cpu_progbuf = n7366; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:131:10  */
  assign dm_ctrl = n7370; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:141:10  */
  assign auth = n7371; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:186:10  */
  assign accen = n7330; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:186:17  */
  assign rden = n7333; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:186:23  */
  assign wren = n7353; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:189:10  */
  assign cpu_rsp_dec = 1'b1; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:202:10  */
  assign dci = n7377; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:209:35  */
  assign n6251 = n6239[8:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:209:38  */
  assign n6253 = n6251 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:209:19  */
  assign n6254 = n6253 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:210:35  */
  assign n6257 = n6239[8:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:210:38  */
  assign n6259 = n6257 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:210:19  */
  assign n6260 = n6259 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:212:29  */
  assign n6263 = 1'b1 ? dmi_wren : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:213:29  */
  assign n6266 = 1'b1 ? dmi_rden : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:220:16  */
  assign n6269 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:229:18  */
  assign n6278 = dm_reg[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:229:37  */
  assign n6279 = ~n6278;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:245:22  */
  assign n6290 = dm_ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:250:29  */
  assign n6291 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:250:34  */
  assign n6293 = n6291 == 7'b0010111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:251:29  */
  assign n6294 = dm_ctrl[41:39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:251:36  */
  assign n6296 = n6294 == 3'b000;
  assign n6298 = dm_ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:250:15  */
  assign n6299 = n6301 ? 3'b001 : n6298;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:250:15  */
  assign n6301 = n6296 & n6293;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:255:27  */
  assign n6302 = dm_reg[113]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:255:57  */
  assign n6303 = dm_reg[112]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:255:46  */
  assign n6304 = n6302 | n6303;
  assign n6306 = dm_ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:255:13  */
  assign n6307 = n6304 ? 3'b001 : n6306;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:249:13  */
  assign n6308 = dmi_wren_auth ? n6299 : n6307;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:247:11  */
  assign n6310 = n6290 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:261:31  */
  assign n6311 = dm_reg[100:93]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:261:46  */
  assign n6313 = n6311 == 8'b00000000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:262:31  */
  assign n6314 = dm_reg[92]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:262:36  */
  assign n6315 = ~n6314;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:261:55  */
  assign n6316 = n6315 & n6313;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:263:31  */
  assign n6317 = dm_reg[91:89]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:263:46  */
  assign n6319 = n6317 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:262:43  */
  assign n6320 = n6319 & n6316;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:264:31  */
  assign n6321 = dm_reg[88]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:264:36  */
  assign n6322 = ~n6321;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:263:55  */
  assign n6323 = n6322 & n6320;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:265:32  */
  assign n6324 = dm_reg[86]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:265:37  */
  assign n6325 = ~n6324;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:265:62  */
  assign n6326 = dm_reg[84:74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:265:76  */
  assign n6328 = n6326 == 11'b00010000000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:265:44  */
  assign n6329 = n6325 | n6328;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:264:43  */
  assign n6330 = n6329 & n6323;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:266:39  */
  assign n6332 = dm_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:266:62  */
  assign n6333 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:266:51  */
  assign n6334 = n6332 & n6333;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6341 = 1'b0 | n6334;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:266:15  */
  assign n6346 = n6341 ? 3'b010 : 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:266:15  */
  assign n6347 = n6341 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:261:13  */
  assign n6350 = n6330 ? n6346 : 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:261:13  */
  assign n6351 = n6330 ? n6347 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:261:13  */
  assign n6352 = n6330 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:259:11  */
  assign n6354 = n6290 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:279:31  */
  assign n6355 = dm_reg[86]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:280:33  */
  assign n6356 = dm_reg[85]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:280:38  */
  assign n6357 = ~n6356;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:283:69  */
  assign n6360 = dm_reg[73:69]; // extract
  assign n6363 = n6281[19:12]; // extract
  assign n6364 = n6281[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:288:69  */
  assign n6368 = dm_reg[73:69]; // extract
  assign n6369 = n6365[19:12]; // extract
  assign n6370 = n6365[6:0]; // extract
  assign n6371 = {12'b111100000000, n6369, n6368, n6370};
  assign n6372 = {7'b1111000, n6360, n6363, 5'b00000, n6364};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:280:15  */
  assign n6373 = n6357 ? n6372 : n6371;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:279:13  */
  assign n6375 = n6355 ? n6373 : 32'b00000000000000000000000000010011;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:293:46  */
  assign n6376 = dm_reg[87]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:277:11  */
  assign n6379 = n6290 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:298:35  */
  assign n6380 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:299:33  */
  assign n6382 = dci[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:299:52  */
  assign n6383 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:299:41  */
  assign n6384 = n6382 & n6383;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6391 = 1'b0 | n6384;
  assign n6394 = dm_ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:299:13  */
  assign n6395 = n6391 ? 3'b100 : n6394;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:296:11  */
  assign n6397 = n6290 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:305:33  */
  assign n6399 = dci[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:305:52  */
  assign n6400 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:305:41  */
  assign n6401 = n6399 & n6400;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6408 = 1'b0 | n6401;
  assign n6411 = dm_ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:305:13  */
  assign n6412 = n6408 ? 3'b000 : n6411;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:303:11  */
  assign n6414 = n6290 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:309:11  */
  assign n6417 = n6290 == 3'b101;
  assign n6419 = {n6417, n6414, n6397, n6379, n6354, n6310};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:245:9  */
  always @*
    case (n6419)
      6'b100000: n6420 = 3'b000;
      6'b010000: n6420 = n6412;
      6'b001000: n6420 = n6395;
      6'b000100: n6420 = 3'b011;
      6'b000010: n6420 = n6350;
      6'b000001: n6420 = n6308;
      default: n6420 = 3'b000;
    endcase
  assign n6421 = dm_ctrl[35:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:245:9  */
  always @*
    case (n6419)
      6'b100000: n6422 = n6421;
      6'b010000: n6422 = n6421;
      6'b001000: n6422 = n6421;
      6'b000100: n6422 = n6375;
      6'b000010: n6422 = n6421;
      6'b000001: n6422 = n6421;
      default: n6422 = n6421;
    endcase
  assign n6423 = dm_ctrl[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:245:9  */
  always @*
    case (n6419)
      6'b100000: n6424 = n6423;
      6'b010000: n6424 = n6423;
      6'b001000: n6424 = n6423;
      6'b000100: n6424 = n6376;
      6'b000010: n6424 = n6423;
      6'b000001: n6424 = n6423;
      default: n6424 = n6423;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:245:9  */
  always @*
    case (n6419)
      6'b100000: n6425 = 1'b0;
      6'b010000: n6425 = 1'b0;
      6'b001000: n6425 = 1'b0;
      6'b000100: n6425 = 1'b0;
      6'b000010: n6425 = n6351;
      6'b000001: n6425 = 1'b0;
      default: n6425 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:245:9  */
  always @*
    case (n6419)
      6'b100000: n6426 = 1'b0;
      6'b010000: n6426 = 1'b0;
      6'b001000: n6426 = 1'b0;
      6'b000100: n6426 = 1'b0;
      6'b000010: n6426 = n6352;
      6'b000001: n6426 = 1'b0;
      default: n6426 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:245:9  */
  always @*
    case (n6419)
      6'b100000: n6427 = 1'b0;
      6'b010000: n6427 = 1'b0;
      6'b001000: n6427 = n6380;
      6'b000100: n6427 = 1'b0;
      6'b000010: n6427 = 1'b0;
      6'b000001: n6427 = 1'b0;
      default: n6427 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:320:21  */
  assign n6428 = dm_ctrl[41:39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:320:28  */
  assign n6430 = n6428 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:321:23  */
  assign n6431 = dm_ctrl[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:323:22  */
  assign n6433 = dci[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:325:26  */
  assign n6435 = dm_ctrl[38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:327:25  */
  assign n6437 = dm_reg[110]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:327:54  */
  assign n6438 = dm_reg[109]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:327:43  */
  assign n6439 = n6437 | n6438;
  assign n6441 = dm_ctrl[41:39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:327:11  */
  assign n6442 = n6439 ? 3'b001 : n6441;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:325:11  */
  assign n6443 = n6435 ? 3'b010 : n6442;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:323:11  */
  assign n6444 = n6433 ? 3'b011 : n6443;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:321:11  */
  assign n6445 = n6431 ? 3'b100 : n6444;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:330:23  */
  assign n6446 = dm_reg[111]; // extract
  assign n6448 = dm_ctrl[41:39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:330:9  */
  assign n6449 = n6446 ? 3'b000 : n6448;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:320:9  */
  assign n6450 = n6430 ? n6445 : n6449;
  assign n6451 = {n6450, n6426, n6425, n6424, n6422};
  assign n6452 = {3'b000, 1'b0, 1'b0, 1'b0, 32'b00000000000000000010000000100011};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:229:7  */
  assign n6453 = n6279 ? 3'b000 : n6420;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:229:7  */
  assign n6454 = n6279 ? n6452 : n6451;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:229:7  */
  assign n6455 = n6279 ? 1'b0 : n6427;
  assign n6462 = {3'b000, 1'b0, 1'b0, 1'b0, 32'b00000000000000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:339:37  */
  assign n6468 = dm_ctrl[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:339:43  */
  assign n6470 = n6468 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:339:23  */
  assign n6471 = n6470 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:346:16  */
  assign n6474 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:355:20  */
  assign n6480 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:357:27  */
  assign n6482 = dci[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:359:27  */
  assign n6484 = dci[2]; // extract
  assign n6486 = dm_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:359:9  */
  assign n6487 = n6484 ? 1'b0 : n6486;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:357:9  */
  assign n6488 = n6482 ? 1'b1 : n6487;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:355:9  */
  assign n6489 = n6480 ? 1'b0 : n6488;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:364:20  */
  assign n6490 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:366:23  */
  assign n6492 = dm_reg[102]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:366:61  */
  assign n6493 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:366:38  */
  assign n6494 = n6493 & n6492;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:368:27  */
  assign n6496 = dci[2]; // extract
  assign n6498 = dm_ctrl[43]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:368:9  */
  assign n6499 = n6496 ? 1'b0 : n6498;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:366:9  */
  assign n6500 = n6494 ? 1'b1 : n6499;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:364:9  */
  assign n6501 = n6490 ? 1'b0 : n6500;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:373:20  */
  assign n6502 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:375:27  */
  assign n6504 = dci[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:377:23  */
  assign n6506 = dm_reg[102]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:377:61  */
  assign n6507 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:377:38  */
  assign n6508 = n6507 & n6506;
  assign n6510 = dm_ctrl[44]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:377:9  */
  assign n6511 = n6508 ? 1'b0 : n6510;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:375:9  */
  assign n6512 = n6504 ? 1'b1 : n6511;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:373:9  */
  assign n6513 = n6502 ? 1'b0 : n6512;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:382:20  */
  assign n6514 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:384:23  */
  assign n6516 = dm_reg[103]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:384:63  */
  assign n6517 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:384:40  */
  assign n6518 = n6517 & n6516;
  assign n6520 = dm_ctrl[45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:384:9  */
  assign n6521 = n6518 ? 1'b0 : n6520;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:382:9  */
  assign n6522 = n6514 ? 1'b1 : n6521;
  assign n6523 = {n6522, n6513, n6501, n6489};
  assign n6526 = {1'b0, 1'b0, 1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:397:16  */
  assign n6530 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:424:21  */
  assign n6550 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:424:26  */
  assign n6552 = n6550 == 7'b0010000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:426:54  */
  assign n6553 = n6239[40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:427:54  */
  assign n6554 = n6239[39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:428:54  */
  assign n6555 = n6239[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:429:54  */
  assign n6556 = n6239[27:25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:430:54  */
  assign n6557 = n6239[10]; // extract
  assign n6558 = {n6556, n6555, n6554, n6553};
  assign n6559 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:425:9  */
  assign n6560 = dmi_wren_auth ? n6557 : n6559;
  assign n6561 = dm_reg[101]; // extract
  assign n6562 = dm_reg[106:104]; // extract
  assign n6563 = {n6562, 1'b0, 1'b0, n6561};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:425:9  */
  assign n6564 = dmi_wren_auth ? n6558 : n6563;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:433:54  */
  assign n6565 = n6239[9]; // extract
  assign n6566 = dm_reg[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:432:9  */
  assign n6567 = dmi_wren ? n6565 : n6566;
  assign n6568 = {n6567, n6560};
  assign n6569 = dm_reg[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:424:7  */
  assign n6570 = n6552 ? n6568 : n6569;
  assign n6571 = dm_reg[101]; // extract
  assign n6572 = dm_reg[106:104]; // extract
  assign n6573 = {n6572, 1'b0, 1'b0, n6571};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:424:7  */
  assign n6574 = n6552 ? n6564 : n6573;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:21  */
  assign n6575 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:26  */
  assign n6577 = n6575 == 7'b0010111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:44  */
  assign n6578 = dmi_wren_auth & n6577;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:83  */
  assign n6579 = dm_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:88  */
  assign n6580 = ~n6579;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:70  */
  assign n6581 = n6580 & n6578;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:108  */
  assign n6582 = dm_ctrl[41:39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:115  */
  assign n6584 = n6582 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:95  */
  assign n6585 = n6584 & n6581;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:439:37  */
  assign n6586 = n6239[40:9]; // extract
  assign n6587 = dm_reg[100:69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:438:7  */
  assign n6588 = n6585 ? n6586 : n6587;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:443:21  */
  assign n6589 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:443:26  */
  assign n6591 = n6589 == 7'b0011000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:443:49  */
  assign n6592 = dmi_wren_auth & n6591;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:443:88  */
  assign n6593 = dm_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:443:93  */
  assign n6594 = ~n6593;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:443:75  */
  assign n6595 = n6594 & n6592;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:444:65  */
  assign n6596 = n6239[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:445:65  */
  assign n6597 = n6239[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:446:65  */
  assign n6598 = n6239[26]; // extract
  assign n6599 = {n6598, n6597, n6596};
  assign n6600 = dm_reg[4:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:443:7  */
  assign n6601 = n6595 ? n6599 : n6600;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:450:22  */
  assign n6602 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:450:27  */
  assign n6604 = n6602 == 7'b0000100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:450:58  */
  assign n6605 = dm_reg[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:450:46  */
  assign n6606 = n6605 & n6604;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:451:22  */
  assign n6607 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:451:27  */
  assign n6609 = n6607 == 7'b0100000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:451:86  */
  assign n6610 = dm_reg[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:451:46  */
  assign n6611 = n6610 & n6609;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:450:92  */
  assign n6612 = n6606 | n6611;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:452:22  */
  assign n6613 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:452:27  */
  assign n6615 = n6613 == 7'b0100001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:452:86  */
  assign n6616 = dm_reg[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:452:46  */
  assign n6617 = n6616 & n6615;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:451:98  */
  assign n6618 = n6612 | n6617;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:450:7  */
  assign n6620 = n6621 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:450:7  */
  assign n6621 = dmi_wren_auth & n6618;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:459:21  */
  assign n6622 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:459:26  */
  assign n6624 = n6622 == 7'b0010110;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:459:47  */
  assign n6625 = dmi_wren_auth & n6624;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:459:92  */
  assign n6626 = n6239[19:17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:459:106  */
  assign n6628 = n6626 == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:459:73  */
  assign n6629 = n6628 & n6625;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:459:7  */
  assign n6631 = n6629 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:464:21  */
  assign n6632 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:464:26  */
  assign n6634 = n6632 == 7'b0100000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:464:45  */
  assign n6635 = dmi_wren_auth & n6634;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:464:84  */
  assign n6636 = dm_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:464:89  */
  assign n6637 = ~n6636;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:464:71  */
  assign n6638 = n6637 & n6635;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:465:40  */
  assign n6639 = n6239[40:9]; // extract
  assign n6640 = dm_reg[68:37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:464:7  */
  assign n6641 = n6638 ? n6639 : n6640;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:469:21  */
  assign n6642 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:469:26  */
  assign n6644 = n6642 == 7'b0100001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:469:45  */
  assign n6645 = dmi_wren_auth & n6644;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:469:84  */
  assign n6646 = dm_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:469:89  */
  assign n6647 = ~n6646;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:469:71  */
  assign n6648 = n6647 & n6645;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:470:40  */
  assign n6649 = n6239[40:9]; // extract
  assign n6650 = dm_reg[36:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:469:7  */
  assign n6651 = n6648 ? n6649 : n6650;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:474:45  */
  assign n6652 = dm_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:474:32  */
  assign n6653 = n6652 & dmi_wren_auth;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:475:22  */
  assign n6654 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:475:27  */
  assign n6656 = n6654 == 7'b0010110;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:475:64  */
  assign n6657 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:475:69  */
  assign n6659 = n6657 == 7'b0010111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:475:50  */
  assign n6660 = n6656 | n6659;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:476:22  */
  assign n6661 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:476:27  */
  assign n6663 = n6661 == 7'b0011000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:475:88  */
  assign n6664 = n6660 | n6663;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:476:64  */
  assign n6665 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:476:69  */
  assign n6667 = n6665 == 7'b0000100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:476:50  */
  assign n6668 = n6664 | n6667;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:477:22  */
  assign n6669 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:477:27  */
  assign n6671 = n6669 == 7'b0100000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:476:88  */
  assign n6672 = n6668 | n6671;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:477:64  */
  assign n6673 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:477:69  */
  assign n6675 = n6673 == 7'b0100001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:477:50  */
  assign n6676 = n6672 | n6675;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:474:57  */
  assign n6677 = n6676 & n6653;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:474:7  */
  assign n6679 = n6677 ? 1'b1 : 1'b0;
  assign n6680 = {n6574, n6588, n6641, n6651, n6601, n6570};
  assign n6681 = {n6620, n6631};
  assign n6688 = {3'b000, 1'b0, 1'b0, 1'b0, 32'b00000000000000000000000000000000, 64'b0000000000000000000000000001001100000000000000000000000000010011, 2'b00, 1'b0, 1'b0, 1'b0};
  assign n6689 = {1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:487:54  */
  assign n6695 = dm_reg[106]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:487:58  */
  assign n6696 = ~n6695;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:487:84  */
  assign n6697 = dm_reg[105:104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:487:97  */
  assign n6699 = n6697 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:487:65  */
  assign n6700 = n6699 & n6696;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:487:34  */
  assign n6701 = n6700 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:489:51  */
  assign n6704 = dm_reg[106:104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:489:60  */
  assign n6706 = $unsigned(n6704) < $unsigned(3'b001);
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:489:29  */
  assign n6707 = n6706 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:495:68  */
  assign n6710 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:495:73  */
  assign n6712 = n6710 == 7'b0000100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:495:53  */
  assign n6713 = n6712 & dmi_wren_auth;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:495:102  */
  assign n6714 = dm_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:495:107  */
  assign n6715 = ~n6714;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:495:89  */
  assign n6716 = n6715 & n6713;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:495:26  */
  assign n6717 = n6716 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:500:30  */
  assign n6719 = dm_reg[101]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:500:61  */
  assign n6720 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:500:39  */
  assign n6721 = n6719 & n6720;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:500:76  */
  assign n6722 = dm_reg[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:500:65  */
  assign n6723 = n6721 & n6722;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:500:95  */
  assign n6725 = 1'b1 ? n6723 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:501:46  */
  assign n6727 = dm_ctrl[43]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:505:33  */
  assign n6729 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:505:71  */
  assign n6730 = dm_reg[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:505:59  */
  assign n6731 = n6730 & n6729;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:505:97  */
  assign n6733 = 1'b1 & n6731;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:505:20  */
  assign n6734 = n6733 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:508:29  */
  assign n6736 = dm_ctrl[35:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:509:47  */
  assign n6737 = dm_ctrl[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:509:55  */
  assign n6738 = ~n6737;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:509:33  */
  assign n6739 = n6738 ? 32'b00000000000000000000000000010011 : n6740;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:509:81  */
  assign n6740 = dm_reg[68:37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:510:47  */
  assign n6741 = dm_ctrl[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:510:55  */
  assign n6742 = ~n6741;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:510:33  */
  assign n6743 = n6742 ? 32'b00000000000000000000000000010011 : n6744;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:510:81  */
  assign n6744 = dm_reg[36:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:518:16  */
  assign n6747 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:524:34  */
  assign n6753 = dmi_wren | dmi_rden;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:22  */
  assign n6755 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:534:65  */
  assign n6760 = dm_ctrl[45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:534:87  */
  assign n6761 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:534:76  */
  assign n6762 = n6760 & n6761;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6769 = 1'b0 | n6762;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:535:65  */
  assign n6772 = dm_ctrl[45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:535:87  */
  assign n6773 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:535:76  */
  assign n6774 = n6772 & n6773;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6781 = 1'b0 | n6774;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:536:65  */
  assign n6784 = dm_ctrl[44]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:536:92  */
  assign n6785 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:536:81  */
  assign n6786 = n6784 & n6785;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6793 = 1'b0 | n6786;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:537:65  */
  assign n6796 = dm_ctrl[44]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:537:92  */
  assign n6797 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:537:81  */
  assign n6798 = n6796 & n6797;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6805 = 1'b0 | n6798;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:538:52  */
  assign n6807 = dm_reg[108]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:539:52  */
  assign n6808 = dm_reg[108]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:540:52  */
  assign n6809 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:541:52  */
  assign n6810 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:542:69  */
  assign n6812 = dm_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:542:92  */
  assign n6813 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:542:81  */
  assign n6814 = n6812 & n6813;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6821 = 1'b0 | n6814;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:542:45  */
  assign n6823 = ~n6821;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:543:69  */
  assign n6825 = dm_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:543:92  */
  assign n6826 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:543:81  */
  assign n6827 = n6825 & n6826;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6834 = 1'b0 | n6827;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:543:45  */
  assign n6836 = ~n6834;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:544:65  */
  assign n6838 = dm_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:544:88  */
  assign n6839 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:544:77  */
  assign n6840 = n6838 & n6839;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6847 = 1'b0 | n6840;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:545:65  */
  assign n6850 = dm_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:545:88  */
  assign n6851 = dm_reg[107]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:545:77  */
  assign n6852 = n6850 & n6851;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n6859 = 1'b0 | n6852;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:549:45  */
  assign n6863 = auth[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:550:45  */
  assign n6864 = auth[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:529:9  */
  assign n6867 = n6755 == 7'b0010001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:562:64  */
  assign n6874 = dm_reg[106:104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:562:55  */
  assign n6876 = {7'b0000000, n6874};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:567:52  */
  assign n6881 = dm_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:569:39  */
  assign n6882 = dm_reg[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:554:9  */
  assign n6884 = n6755 == 7'b0010000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:572:9  */
  assign n6892 = n6755 == 7'b0010010;
  assign n6895 = n6893[7:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:587:53  */
  assign n6896 = dm_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:589:53  */
  assign n6898 = dm_ctrl[41:39]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:583:9  */
  assign n6902 = n6755 == 7'b0010110;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:597:42  */
  assign n6903 = dm_reg[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:598:70  */
  assign n6904 = dm_reg[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:599:70  */
  assign n6905 = dm_reg[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:595:9  */
  assign n6907 = n6755 == 7'b0011000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:605:35  */
  assign n6908 = dci[38:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:603:9  */
  assign n6910 = n6755 == 7'b0000100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:610:34  */
  assign n6911 = auth[35:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:609:9  */
  assign n6913 = n6755 == 7'b0110000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:615:72  */
  assign n6914 = dm_ctrl[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:613:9  */
  assign n6916 = n6755 == 7'b1000000;
  assign n6918 = {n6916, n6913, n6910, n6907, n6902, n6892, n6884, n6867};
  assign n6919 = n6865[0]; // extract
  assign n6920 = n6890[0]; // extract
  assign n6921 = n6900[0]; // extract
  assign n6922 = n6908[0]; // extract
  assign n6923 = n6911[0]; // extract
  assign n6924 = n6917[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6925 = n6914;
      8'b01000000: n6925 = n6923;
      8'b00100000: n6925 = n6922;
      8'b00010000: n6925 = n6903;
      8'b00001000: n6925 = n6921;
      8'b00000100: n6925 = n6920;
      8'b00000010: n6925 = n6882;
      8'b00000001: n6925 = n6919;
      default: n6925 = n6924;
    endcase
  assign n6926 = n6865[1]; // extract
  assign n6927 = n6890[1]; // extract
  assign n6928 = n6900[1]; // extract
  assign n6929 = n6908[1]; // extract
  assign n6930 = n6911[1]; // extract
  assign n6931 = n6917[1]; // extract
  assign n6932 = n6754[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6933 = n6932;
      8'b01000000: n6933 = n6930;
      8'b00100000: n6933 = n6929;
      8'b00010000: n6933 = n6932;
      8'b00001000: n6933 = n6928;
      8'b00000100: n6933 = n6927;
      8'b00000010: n6933 = n6881;
      8'b00000001: n6933 = n6926;
      default: n6933 = n6931;
    endcase
  assign n6934 = n6865[2]; // extract
  assign n6935 = n6890[2]; // extract
  assign n6936 = n6900[2]; // extract
  assign n6937 = n6908[2]; // extract
  assign n6938 = n6911[2]; // extract
  assign n6939 = n6917[2]; // extract
  assign n6940 = n6754[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6941 = n6940;
      8'b01000000: n6941 = n6938;
      8'b00100000: n6941 = n6937;
      8'b00010000: n6941 = n6940;
      8'b00001000: n6941 = n6936;
      8'b00000100: n6941 = n6935;
      8'b00000010: n6941 = 1'b0;
      8'b00000001: n6941 = n6934;
      default: n6941 = n6939;
    endcase
  assign n6942 = n6865[3]; // extract
  assign n6943 = n6890[3]; // extract
  assign n6944 = n6900[3]; // extract
  assign n6945 = n6908[3]; // extract
  assign n6946 = n6911[3]; // extract
  assign n6947 = n6917[3]; // extract
  assign n6948 = n6754[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6949 = n6948;
      8'b01000000: n6949 = n6946;
      8'b00100000: n6949 = n6945;
      8'b00010000: n6949 = n6948;
      8'b00001000: n6949 = n6944;
      8'b00000100: n6949 = n6943;
      8'b00000010: n6949 = 1'b0;
      8'b00000001: n6949 = n6942;
      default: n6949 = n6947;
    endcase
  assign n6950 = n6878[0]; // extract
  assign n6951 = n6890[4]; // extract
  assign n6952 = n6899[0]; // extract
  assign n6953 = n6908[4]; // extract
  assign n6954 = n6911[4]; // extract
  assign n6955 = n6917[4]; // extract
  assign n6956 = n6754[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6957 = n6956;
      8'b01000000: n6957 = n6954;
      8'b00100000: n6957 = n6953;
      8'b00010000: n6957 = n6956;
      8'b00001000: n6957 = n6952;
      8'b00000100: n6957 = n6951;
      8'b00000010: n6957 = n6950;
      8'b00000001: n6957 = 1'b0;
      default: n6957 = n6955;
    endcase
  assign n6958 = n6878[1]; // extract
  assign n6959 = n6890[5]; // extract
  assign n6960 = n6899[1]; // extract
  assign n6961 = n6908[5]; // extract
  assign n6962 = n6911[5]; // extract
  assign n6963 = n6917[5]; // extract
  assign n6964 = n6754[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6965 = n6964;
      8'b01000000: n6965 = n6962;
      8'b00100000: n6965 = n6961;
      8'b00010000: n6965 = n6964;
      8'b00001000: n6965 = n6960;
      8'b00000100: n6965 = n6959;
      8'b00000010: n6965 = n6958;
      8'b00000001: n6965 = 1'b0;
      default: n6965 = n6963;
    endcase
  assign n6966 = n6877[0]; // extract
  assign n6967 = n6890[6]; // extract
  assign n6968 = n6899[2]; // extract
  assign n6969 = n6908[6]; // extract
  assign n6970 = n6911[6]; // extract
  assign n6971 = n6917[6]; // extract
  assign n6972 = n6754[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6973 = n6972;
      8'b01000000: n6973 = n6970;
      8'b00100000: n6973 = n6969;
      8'b00010000: n6973 = n6972;
      8'b00001000: n6973 = n6968;
      8'b00000100: n6973 = n6967;
      8'b00000010: n6973 = n6966;
      8'b00000001: n6973 = n6864;
      default: n6973 = n6971;
    endcase
  assign n6974 = n6877[1]; // extract
  assign n6975 = n6890[7]; // extract
  assign n6976 = n6899[3]; // extract
  assign n6977 = n6908[7]; // extract
  assign n6978 = n6911[7]; // extract
  assign n6979 = n6917[7]; // extract
  assign n6980 = n6754[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6981 = n6980;
      8'b01000000: n6981 = n6978;
      8'b00100000: n6981 = n6977;
      8'b00010000: n6981 = n6980;
      8'b00001000: n6981 = n6976;
      8'b00000100: n6981 = n6975;
      8'b00000010: n6981 = n6974;
      8'b00000001: n6981 = n6863;
      default: n6981 = n6979;
    endcase
  assign n6982 = n6877[2]; // extract
  assign n6983 = n6890[8]; // extract
  assign n6984 = n6898[0]; // extract
  assign n6985 = n6908[8]; // extract
  assign n6986 = n6911[8]; // extract
  assign n6987 = n6917[8]; // extract
  assign n6988 = n6754[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6989 = n6988;
      8'b01000000: n6989 = n6986;
      8'b00100000: n6989 = n6985;
      8'b00010000: n6989 = n6988;
      8'b00001000: n6989 = n6984;
      8'b00000100: n6989 = n6983;
      8'b00000010: n6989 = n6982;
      8'b00000001: n6989 = n6859;
      default: n6989 = n6987;
    endcase
  assign n6990 = n6877[3]; // extract
  assign n6991 = n6890[9]; // extract
  assign n6992 = n6898[1]; // extract
  assign n6993 = n6908[9]; // extract
  assign n6994 = n6911[9]; // extract
  assign n6995 = n6917[9]; // extract
  assign n6996 = n6754[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n6997 = n6996;
      8'b01000000: n6997 = n6994;
      8'b00100000: n6997 = n6993;
      8'b00010000: n6997 = n6996;
      8'b00001000: n6997 = n6992;
      8'b00000100: n6997 = n6991;
      8'b00000010: n6997 = n6990;
      8'b00000001: n6997 = n6847;
      default: n6997 = n6995;
    endcase
  assign n6998 = n6877[4]; // extract
  assign n6999 = n6890[10]; // extract
  assign n7000 = n6898[2]; // extract
  assign n7001 = n6908[10]; // extract
  assign n7002 = n6911[10]; // extract
  assign n7003 = n6917[10]; // extract
  assign n7004 = n6754[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7005 = n7004;
      8'b01000000: n7005 = n7002;
      8'b00100000: n7005 = n7001;
      8'b00010000: n7005 = n7004;
      8'b00001000: n7005 = n7000;
      8'b00000100: n7005 = n6999;
      8'b00000010: n7005 = n6998;
      8'b00000001: n7005 = n6836;
      default: n7005 = n7003;
    endcase
  assign n7006 = n6877[5]; // extract
  assign n7007 = n6890[11]; // extract
  assign n7008 = n6908[11]; // extract
  assign n7009 = n6911[11]; // extract
  assign n7010 = n6917[11]; // extract
  assign n7011 = n6754[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7012 = n7011;
      8'b01000000: n7012 = n7009;
      8'b00100000: n7012 = n7008;
      8'b00010000: n7012 = n7011;
      8'b00001000: n7012 = 1'b1;
      8'b00000100: n7012 = n7007;
      8'b00000010: n7012 = n7006;
      8'b00000001: n7012 = n6823;
      default: n7012 = n7010;
    endcase
  assign n7013 = n6877[6]; // extract
  assign n7014 = n6889[0]; // extract
  assign n7015 = n6908[12]; // extract
  assign n7016 = n6911[12]; // extract
  assign n7017 = n6917[12]; // extract
  assign n7018 = n6754[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7019 = n7018;
      8'b01000000: n7019 = n7016;
      8'b00100000: n7019 = n7015;
      8'b00010000: n7019 = n7018;
      8'b00001000: n7019 = n6896;
      8'b00000100: n7019 = n7014;
      8'b00000010: n7019 = n7013;
      8'b00000001: n7019 = n6810;
      default: n7019 = n7017;
    endcase
  assign n7020 = n6877[7]; // extract
  assign n7021 = n6889[1]; // extract
  assign n7022 = n6908[13]; // extract
  assign n7023 = n6911[13]; // extract
  assign n7024 = n6917[13]; // extract
  assign n7025 = n6754[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7026 = n7025;
      8'b01000000: n7026 = n7023;
      8'b00100000: n7026 = n7022;
      8'b00010000: n7026 = n7025;
      8'b00001000: n7026 = n7025;
      8'b00000100: n7026 = n7021;
      8'b00000010: n7026 = n7020;
      8'b00000001: n7026 = n6809;
      default: n7026 = n7024;
    endcase
  assign n7027 = n6877[8]; // extract
  assign n7028 = n6889[2]; // extract
  assign n7029 = n6908[14]; // extract
  assign n7030 = n6911[14]; // extract
  assign n7031 = n6917[14]; // extract
  assign n7032 = n6754[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7033 = n7032;
      8'b01000000: n7033 = n7030;
      8'b00100000: n7033 = n7029;
      8'b00010000: n7033 = n7032;
      8'b00001000: n7033 = n7032;
      8'b00000100: n7033 = n7028;
      8'b00000010: n7033 = n7027;
      8'b00000001: n7033 = n6808;
      default: n7033 = n7031;
    endcase
  assign n7034 = n6877[9]; // extract
  assign n7035 = n6889[3]; // extract
  assign n7036 = n6908[15]; // extract
  assign n7037 = n6911[15]; // extract
  assign n7038 = n6917[15]; // extract
  assign n7039 = n6754[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7040 = n7039;
      8'b01000000: n7040 = n7037;
      8'b00100000: n7040 = n7036;
      8'b00010000: n7040 = n7039;
      8'b00001000: n7040 = n7039;
      8'b00000100: n7040 = n7035;
      8'b00000010: n7040 = n7034;
      8'b00000001: n7040 = n6807;
      default: n7040 = n7038;
    endcase
  assign n7041 = n6876[0]; // extract
  assign n7042 = n6908[16]; // extract
  assign n7043 = n6911[16]; // extract
  assign n7044 = n6917[16]; // extract
  assign n7045 = n6754[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7046 = n7045;
      8'b01000000: n7046 = n7043;
      8'b00100000: n7046 = n7042;
      8'b00010000: n7046 = n6904;
      8'b00001000: n7046 = n7045;
      8'b00000100: n7046 = 1'b1;
      8'b00000010: n7046 = n7041;
      8'b00000001: n7046 = n6805;
      default: n7046 = n7044;
    endcase
  assign n7047 = n6876[1]; // extract
  assign n7048 = n6887[0]; // extract
  assign n7049 = n6908[17]; // extract
  assign n7050 = n6911[17]; // extract
  assign n7051 = n6917[17]; // extract
  assign n7052 = n6754[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7053 = n7052;
      8'b01000000: n7053 = n7050;
      8'b00100000: n7053 = n7049;
      8'b00010000: n7053 = n6905;
      8'b00001000: n7053 = n7052;
      8'b00000100: n7053 = n7048;
      8'b00000010: n7053 = n7047;
      8'b00000001: n7053 = n6793;
      default: n7053 = n7051;
    endcase
  assign n7054 = n6876[2]; // extract
  assign n7055 = n6887[1]; // extract
  assign n7056 = n6908[18]; // extract
  assign n7057 = n6911[18]; // extract
  assign n7058 = n6917[18]; // extract
  assign n7059 = n6754[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7060 = n7059;
      8'b01000000: n7060 = n7057;
      8'b00100000: n7060 = n7056;
      8'b00010000: n7060 = n7059;
      8'b00001000: n7060 = n7059;
      8'b00000100: n7060 = n7055;
      8'b00000010: n7060 = n7054;
      8'b00000001: n7060 = n6781;
      default: n7060 = n7058;
    endcase
  assign n7061 = n6876[3]; // extract
  assign n7062 = n6887[2]; // extract
  assign n7063 = n6908[19]; // extract
  assign n7064 = n6911[19]; // extract
  assign n7065 = n6917[19]; // extract
  assign n7066 = n6754[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7067 = n7066;
      8'b01000000: n7067 = n7064;
      8'b00100000: n7067 = n7063;
      8'b00010000: n7067 = n7066;
      8'b00001000: n7067 = n7066;
      8'b00000100: n7067 = n7062;
      8'b00000010: n7067 = n7061;
      8'b00000001: n7067 = n6769;
      default: n7067 = n7065;
    endcase
  assign n7068 = n6876[5:4]; // extract
  assign n7069 = n6886[1:0]; // extract
  assign n7070 = n6908[21:20]; // extract
  assign n7071 = n6911[21:20]; // extract
  assign n7072 = n6917[21:20]; // extract
  assign n7073 = n6754[21:20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7074 = n7073;
      8'b01000000: n7074 = n7071;
      8'b00100000: n7074 = n7070;
      8'b00010000: n7074 = n7073;
      8'b00001000: n7074 = n7073;
      8'b00000100: n7074 = n7069;
      8'b00000010: n7074 = n7068;
      8'b00000001: n7074 = 2'b00;
      default: n7074 = n7072;
    endcase
  assign n7075 = n6876[6]; // extract
  assign n7076 = n6886[2]; // extract
  assign n7077 = n6908[22]; // extract
  assign n7078 = n6911[22]; // extract
  assign n7079 = n6917[22]; // extract
  assign n7080 = n6754[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7081 = n7080;
      8'b01000000: n7081 = n7078;
      8'b00100000: n7081 = n7077;
      8'b00010000: n7081 = n7080;
      8'b00001000: n7081 = n7080;
      8'b00000100: n7081 = n7076;
      8'b00000010: n7081 = n7075;
      8'b00000001: n7081 = 1'b1;
      default: n7081 = n7079;
    endcase
  assign n7082 = n6756[0]; // extract
  assign n7083 = n6876[7]; // extract
  assign n7084 = n6886[3]; // extract
  assign n7085 = n6908[23]; // extract
  assign n7086 = n6911[23]; // extract
  assign n7087 = n6917[23]; // extract
  assign n7088 = n6754[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7089 = n7088;
      8'b01000000: n7089 = n7086;
      8'b00100000: n7089 = n7085;
      8'b00010000: n7089 = n7088;
      8'b00001000: n7089 = n7088;
      8'b00000100: n7089 = n7084;
      8'b00000010: n7089 = n7083;
      8'b00000001: n7089 = n7082;
      default: n7089 = n7087;
    endcase
  assign n7090 = n6756[2:1]; // extract
  assign n7091 = n6876[9:8]; // extract
  assign n7092 = n6885[1:0]; // extract
  assign n7093 = n6894[1:0]; // extract
  assign n7094 = n6908[25:24]; // extract
  assign n7095 = n6911[25:24]; // extract
  assign n7096 = n6917[25:24]; // extract
  assign n7097 = n6754[25:24]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7098 = n7097;
      8'b01000000: n7098 = n7095;
      8'b00100000: n7098 = n7094;
      8'b00010000: n7098 = n7097;
      8'b00001000: n7098 = n7093;
      8'b00000100: n7098 = n7092;
      8'b00000010: n7098 = n7091;
      8'b00000001: n7098 = n7090;
      default: n7098 = n7096;
    endcase
  assign n7099 = n6756[3]; // extract
  assign n7100 = n6885[2]; // extract
  assign n7101 = n6894[2]; // extract
  assign n7102 = n6908[26]; // extract
  assign n7103 = n6911[26]; // extract
  assign n7104 = n6917[26]; // extract
  assign n7105 = n6754[26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7106 = n7105;
      8'b01000000: n7106 = n7103;
      8'b00100000: n7106 = n7102;
      8'b00010000: n7106 = n7105;
      8'b00001000: n7106 = n7101;
      8'b00000100: n7106 = n7100;
      8'b00000010: n7106 = 1'b0;
      8'b00000001: n7106 = n7099;
      default: n7106 = n7104;
    endcase
  assign n7107 = n6756[4]; // extract
  assign n7108 = n6885[3]; // extract
  assign n7109 = n6894[3]; // extract
  assign n7110 = n6908[27]; // extract
  assign n7111 = n6911[27]; // extract
  assign n7112 = n6917[27]; // extract
  assign n7113 = n6754[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7114 = n7113;
      8'b01000000: n7114 = n7111;
      8'b00100000: n7114 = n7110;
      8'b00010000: n7114 = n7113;
      8'b00001000: n7114 = n7109;
      8'b00000100: n7114 = n7108;
      8'b00000010: n7114 = 1'b0;
      8'b00000001: n7114 = n7107;
      default: n7114 = n7112;
    endcase
  assign n7115 = n6756[5]; // extract
  assign n7116 = n6885[4]; // extract
  assign n7117 = n6894[4]; // extract
  assign n7118 = n6908[28]; // extract
  assign n7119 = n6911[28]; // extract
  assign n7120 = n6917[28]; // extract
  assign n7121 = n6754[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7122 = n7121;
      8'b01000000: n7122 = n7119;
      8'b00100000: n7122 = n7118;
      8'b00010000: n7122 = n7121;
      8'b00001000: n7122 = n7117;
      8'b00000100: n7122 = n7116;
      8'b00000010: n7122 = 1'b0;
      8'b00000001: n7122 = n7115;
      default: n7122 = n7120;
    endcase
  assign n7123 = n6756[6]; // extract
  assign n7124 = n6885[5]; // extract
  assign n7125 = n6895[0]; // extract
  assign n7126 = n6908[29]; // extract
  assign n7127 = n6911[29]; // extract
  assign n7128 = n6917[29]; // extract
  assign n7129 = n6754[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7130 = n7129;
      8'b01000000: n7130 = n7127;
      8'b00100000: n7130 = n7126;
      8'b00010000: n7130 = n7129;
      8'b00001000: n7130 = n7125;
      8'b00000100: n7130 = n7124;
      8'b00000010: n7130 = 1'b0;
      8'b00000001: n7130 = n7123;
      default: n7130 = n7128;
    endcase
  assign n7131 = n6756[7]; // extract
  assign n7132 = n6885[6]; // extract
  assign n7133 = n6895[1]; // extract
  assign n7134 = n6908[30]; // extract
  assign n7135 = n6911[30]; // extract
  assign n7136 = n6917[30]; // extract
  assign n7137 = n6754[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7138 = n7137;
      8'b01000000: n7138 = n7135;
      8'b00100000: n7138 = n7134;
      8'b00010000: n7138 = n7137;
      8'b00001000: n7138 = n7133;
      8'b00000100: n7138 = n7132;
      8'b00000010: n7138 = 1'b0;
      8'b00000001: n7138 = n7131;
      default: n7138 = n7136;
    endcase
  assign n7139 = n6756[8]; // extract
  assign n7140 = n6885[7]; // extract
  assign n7141 = n6895[2]; // extract
  assign n7142 = n6908[31]; // extract
  assign n7143 = n6911[31]; // extract
  assign n7144 = n6917[31]; // extract
  assign n7145 = n6754[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:526:7  */
  always @*
    case (n6918)
      8'b10000000: n7146 = n7145;
      8'b01000000: n7146 = n7143;
      8'b00100000: n7146 = n7142;
      8'b00010000: n7146 = n7145;
      8'b00001000: n7146 = n7141;
      8'b00000100: n7146 = n7140;
      8'b00000010: n7146 = 1'b0;
      8'b00000001: n7146 = n7139;
      default: n7146 = n7144;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:626:45  */
  assign n7176 = dm_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:626:32  */
  assign n7177 = n7176 & dmi_rden_auth;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:627:22  */
  assign n7178 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:627:27  */
  assign n7180 = n7178 == 7'b0000100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:627:57  */
  assign n7181 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:627:62  */
  assign n7183 = n7181 == 7'b0100000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:627:43  */
  assign n7184 = n7180 | n7183;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:627:95  */
  assign n7185 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:627:100  */
  assign n7187 = n7185 == 7'b0100001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:627:81  */
  assign n7188 = n7184 | n7187;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:626:57  */
  assign n7189 = n7188 & n7177;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:626:7  */
  assign n7192 = n7189 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:636:23  */
  assign n7193 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:636:28  */
  assign n7195 = n7193 == 7'b0000100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:636:59  */
  assign n7196 = dm_reg[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:636:47  */
  assign n7197 = n7196 & n7195;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:637:23  */
  assign n7198 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:637:28  */
  assign n7200 = n7198 == 7'b0100000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:637:87  */
  assign n7201 = dm_reg[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:637:47  */
  assign n7202 = n7201 & n7200;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:636:99  */
  assign n7203 = n7197 | n7202;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:638:23  */
  assign n7204 = n6239[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:638:28  */
  assign n7206 = n7204 == 7'b0100001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:638:87  */
  assign n7207 = dm_reg[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:638:47  */
  assign n7208 = n7207 & n7206;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:637:99  */
  assign n7209 = n7203 | n7208;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:635:32  */
  assign n7210 = n7209 & dmi_rden_auth;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:635:7  */
  assign n7213 = n7210 ? 1'b1 : 1'b0;
  assign n7214 = {n6753, n7146, n7138, n7130, n7122, n7114, n7106, n7098, n7089, n7081, n7074, n7067, n7060, n7053, n7046, n7040, n7033, n7026, n7019, n7012, n7005, n6997, n6989, n6981, n6973, n6965, n6957, n6949, n6941, n6933, n6925};
  assign n7220 = {1'b0, 32'b00000000000000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:652:16  */
  assign n7226 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:665:15  */
  assign n7234 = dci[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:666:35  */
  assign n7235 = n6239[40:9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:667:45  */
  assign n7236 = n6243[8:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:667:58  */
  assign n7238 = n7236 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:667:26  */
  assign n7239 = n7238 & wren;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:668:35  */
  assign n7240 = n6243[63:32]; // extract
  assign n7241 = dci[38:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:667:7  */
  assign n7242 = n7239 ? n7240 : n7241;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:665:7  */
  assign n7243 = n7234 ? n7235 : n7242;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:676:42  */
  assign n7248 = n6243[8:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:676:55  */
  assign n7250 = n7248 == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:676:23  */
  assign n7251 = n7250 & wren;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:678:30  */
  assign n7252 = n6243[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:679:13  */
  assign n7254 = n7252 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:680:13  */
  assign n7256 = n7252 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:681:13  */
  assign n7258 = n7252 == 2'b10;
  assign n7260 = {n7258, n7256, n7254};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:678:11  */
  always @*
    case (n7260)
      3'b100: n7261 = 1'b0;
      3'b010: n7261 = 1'b0;
      3'b001: n7261 = cpu_rsp_dec;
      default: n7261 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:678:11  */
  always @*
    case (n7260)
      3'b100: n7262 = 1'b0;
      3'b010: n7262 = cpu_rsp_dec;
      3'b001: n7262 = 1'b0;
      default: n7262 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:678:11  */
  always @*
    case (n7260)
      3'b100: n7263 = cpu_rsp_dec;
      3'b010: n7263 = 1'b0;
      3'b001: n7263 = 1'b0;
      default: n7263 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:678:11  */
  always @*
    case (n7260)
      3'b100: n7264 = 1'b0;
      3'b010: n7264 = 1'b0;
      3'b001: n7264 = 1'b0;
      default: n7264 = 1'b1;
    endcase
  assign n7265 = {n7264, n7263};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:676:7  */
  assign n7266 = n7251 ? n7261 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:676:7  */
  assign n7267 = n7251 ? n7262 : 1'b0;
  assign n7268 = {1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:676:7  */
  assign n7269 = n7251 ? n7265 : n7268;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:690:28  */
  assign n7271 = n6243[8:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:692:76  */
  assign n7272 = n6243[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:691:11  */
  assign n7280 = n7271 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:694:77  */
  assign n7281 = n6243[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:694:43  */
  assign n7284 = 2'b11 - n7281;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:693:11  */
  assign n7288 = n7271 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:696:35  */
  assign n7289 = dci[38:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:695:11  */
  assign n7291 = n7271 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:699:51  */
  assign n7292 = dci[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:700:51  */
  assign n7293 = dci[3]; // extract
  assign n7294 = {n7291, n7288, n7280};
  assign n7295 = n7382[0]; // extract
  assign n7296 = n7383[0]; // extract
  assign n7297 = n7289[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:690:9  */
  always @*
    case (n7294)
      3'b100: n7298 = n7297;
      3'b010: n7298 = n7296;
      3'b001: n7298 = n7295;
      default: n7298 = n7292;
    endcase
  assign n7299 = n7382[1]; // extract
  assign n7300 = n7383[1]; // extract
  assign n7301 = n7289[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:690:9  */
  always @*
    case (n7294)
      3'b100: n7302 = n7301;
      3'b010: n7302 = n7300;
      3'b001: n7302 = n7299;
      default: n7302 = n7293;
    endcase
  assign n7303 = n7382[31:2]; // extract
  assign n7304 = n7383[31:2]; // extract
  assign n7305 = n7289[31:2]; // extract
  assign n7306 = n7270[31:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:690:9  */
  always @*
    case (n7294)
      3'b100: n7307 = n7305;
      3'b010: n7307 = n7304;
      3'b001: n7307 = n7303;
      default: n7307 = n7306;
    endcase
  assign n7308 = {n7307, n7302, n7298};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:689:7  */
  assign n7309 = rden ? n7308 : 32'b00000000000000000000000000000000;
  assign n7310 = {1'b0, accen, n7309};
  assign n7322 = {1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:708:22  */
  assign n7328 = n6243[79]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:708:42  */
  assign n7329 = n6243[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:708:28  */
  assign n7330 = n7328 & n7329;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:709:37  */
  assign n7331 = n6243[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:709:23  */
  assign n7332 = ~n7331;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:709:18  */
  assign n7333 = accen & n7332;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:710:37  */
  assign n7334 = n6243[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:710:18  */
  assign n7335 = accen & n7334;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n7343 = n6243[67]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n7345 = 1'b1 & n7343;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n7347 = n6243[66]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n7348 = n7345 & n7347;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n7349 = n6243[65]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n7350 = n7348 & n7349;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n7351 = n6243[64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n7352 = n7350 & n7351;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:710:41  */
  assign n7353 = n7335 & n7352;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:523:5  */
  always @(posedge clk_i or posedge n6747)
    if (n6747)
      n7360 <= 1'b0;
    else
      n7360 <= n7213;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:523:5  */
  always @(posedge clk_i or posedge n6747)
    if (n6747)
      n7361 <= 1'b0;
    else
      n7361 <= n7192;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:414:5  */
  always @(posedge clk_i or posedge n6530)
    if (n6530)
      n7362 <= n6689;
    else
      n7362 <= n6681;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:414:5  */
  always @(posedge clk_i or posedge n6530)
    if (n6530)
      n7363 <= 1'b0;
    else
      n7363 <= n6679;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:414:5  */
  always @(posedge clk_i or posedge n6530)
    if (n6530)
      n7364 <= n6688;
    else
      n7364 <= n6680;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:397:5  */
  assign n7365 = {n7360, n7362, n7361, n7363, n6707, n6701, n7364};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:397:5  */
  assign n7366 = {n6736, n6739, n6743, 32'b00000000000100000000000001110011};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:351:5  */
  always @(posedge clk_i or posedge n6474)
    if (n6474)
      n7367 <= n6526;
    else
      n7367 <= n6523;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:228:5  */
  always @(posedge clk_i or posedge n6269)
    if (n6269)
      n7368 <= n6462;
    else
      n7368 <= n6454;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:228:5  */
  always @(posedge clk_i or posedge n6269)
    if (n6269)
      n7369 <= 3'b000;
    else
      n7369 <= n6453;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:220:5  */
  assign n7370 = {n7367, n7368, n6471, n7369};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:220:5  */
  assign n7371 = {32'b00000000000000000000000000000000, 1'b0, 1'b0, 1'b1, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:659:5  */
  always @(posedge clk_i or posedge n7226)
    if (n7226)
      n7372 <= 32'b00000000000000000000000000000000;
    else
      n7372 <= n7243;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:659:5  */
  always @(posedge clk_i or posedge n7226)
    if (n7226)
      n7373 <= n7322;
    else
      n7373 <= n7269;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:659:5  */
  always @(posedge clk_i or posedge n7226)
    if (n7226)
      n7374 <= 1'b0;
    else
      n7374 <= n7267;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:659:5  */
  always @(posedge clk_i or posedge n7226)
    if (n7226)
      n7375 <= 1'b0;
    else
      n7375 <= n7266;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:228:5  */
  always @(posedge clk_i or posedge n6269)
    if (n6269)
      n7376 <= 1'b0;
    else
      n7376 <= n6455;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:220:5  */
  assign n7377 = {n7372, n6717, n7373, n7376, n7374, n6727, n7375};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:523:5  */
  always @(posedge clk_i or posedge n6747)
    if (n6747)
      n7378 <= n7220;
    else
      n7378 <= n7214;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:659:5  */
  always @(posedge clk_i or posedge n7226)
    if (n7226)
      n7379 <= 34'b0000000000000000000000000000000000;
    else
      n7379 <= n7310;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:692:42  */
  reg [31:0] n7380[31:0] ; // memory
  initial begin
    n7380[31] = 32'b00000000000000000000000001110011;
    n7380[30] = 32'b00000000000000000000000001110011;
    n7380[29] = 32'b00000000000000000000000001110011;
    n7380[28] = 32'b00000000000000000000000001110011;
    n7380[27] = 32'b00000000000000000000000001110011;
    n7380[26] = 32'b00000000000000000000000001110011;
    n7380[25] = 32'b00000000000000000000000001110011;
    n7380[24] = 32'b00000000000000000000000001110011;
    n7380[23] = 32'b11101000000000000000000001100111;
    n7380[22] = 32'b00000000000000000001000000001111;
    n7380[21] = 32'b01111011001000000010010001110011;
    n7380[20] = 32'b11111000100000000010010000100011;
    n7380[19] = 32'b11110001010000000010010001110011;
    n7380[18] = 32'b01111011001000000000000001110011;
    n7380[17] = 32'b01111011001000000010010001110011;
    n7380[16] = 32'b11111000100000000010001000100011;
    n7380[15] = 32'b11110001010000000010010001110011;
    n7380[14] = 32'b11111110000001000000001011100011;
    n7380[13] = 32'b00000000000101000111010000010011;
    n7380[12] = 32'b11111000000001000100010000000011;
    n7380[11] = 32'b11110001010000000010010001110011;
    n7380[10] = 32'b00000010000001000001001001100011;
    n7380[9] = 32'b00000000001001000111010000010011;
    n7380[8] = 32'b11111000000001000100010000000011;
    n7380[7] = 32'b11110001010000000010010001110011;
    n7380[6] = 32'b11111000100000000010000000100011;
    n7380[5] = 32'b11110001010000000010010001110011;
    n7380[4] = 32'b01111011001001000001000001110011;
    n7380[3] = 32'b00000000000000000000000000010011;
    n7380[2] = 32'b00000000000100000000000001110011;
    n7380[1] = 32'b01111011001000000010010001110011;
    n7380[0] = 32'b11111000000000000010011000100011;
    end
  assign n7382 = n7380[n7272];
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:692:42  */
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dm.vhd:694:43  */
  assign n7383 = cpu_progbuf[n7284 * 32 +: 32]; //(Bmux)
endmodule

module neorv32_debug_dtm_46d1c9a201904415cbd5c7cc672d1649ed497f22
  (input  clk_i,
   input  rstn_i,
   input  jtag_tck_i,
   input  jtag_tdi_i,
   input  jtag_tms_i,
   input  [31:0] \dmi_rsp_i_dmi_rsp_i[data] ,
   input  \dmi_rsp_i_dmi_rsp_i[ack] ,
   input  jtagspi_sdi_i,
   output jtag_tdo_o,
   output [6:0] \dmi_req_o_dmi_req_o[addr] ,
   output [1:0] \dmi_req_o_dmi_req_o[op] ,
   output [31:0] \dmi_req_o_dmi_req_o[data] ,
   output jtagspi_sck_o,
   output jtagspi_sdo_o,
   output jtagspi_csn_o);
  wire [6:0] n5767;
  wire [1:0] n5768;
  wire [31:0] n5769;
  wire [32:0] n5770;
  wire [13:0] tap_sync;
  wire [3:0] tap_ctrl_state;
  wire [185:0] tap_reg;
  wire [2:0] dr_trigger;
  wire [76:0] dmi_ctrl;
  wire n5775;
  wire [1:0] n5780;
  wire [2:0] n5781;
  wire [1:0] n5782;
  wire [2:0] n5783;
  wire [1:0] n5784;
  wire [2:0] n5785;
  wire [8:0] n5786;
  wire [8:0] n5789;
  wire [1:0] n5793;
  wire n5795;
  wire n5796;
  wire [1:0] n5799;
  wire n5801;
  wire n5802;
  wire n5804;
  wire n5805;
  wire n5806;
  wire n5807;
  wire n5808;
  wire n5809;
  wire n5810;
  wire n5811;
  wire n5812;
  wire n5814;
  wire n5816;
  wire n5817;
  wire n5818;
  wire [3:0] n5821;
  wire n5823;
  wire n5824;
  wire n5825;
  wire [3:0] n5828;
  wire n5830;
  wire n5831;
  wire n5832;
  wire [3:0] n5835;
  wire n5837;
  wire n5838;
  wire n5839;
  wire [3:0] n5842;
  wire n5844;
  wire n5845;
  wire n5846;
  wire [3:0] n5849;
  wire n5851;
  wire n5852;
  wire n5853;
  wire [3:0] n5856;
  wire n5858;
  wire n5859;
  wire n5860;
  wire [3:0] n5863;
  wire n5865;
  wire n5866;
  wire n5867;
  wire [3:0] n5870;
  wire n5872;
  wire n5873;
  wire n5874;
  wire [3:0] n5877;
  wire n5879;
  wire n5880;
  wire n5881;
  wire [3:0] n5884;
  wire n5886;
  wire n5887;
  wire n5888;
  wire [3:0] n5891;
  wire n5893;
  wire n5894;
  wire n5895;
  wire [3:0] n5898;
  wire n5900;
  wire n5901;
  wire n5902;
  wire [3:0] n5905;
  wire n5907;
  wire n5908;
  wire n5909;
  wire [3:0] n5912;
  wire n5914;
  wire n5915;
  wire n5916;
  wire [3:0] n5919;
  wire n5921;
  wire n5922;
  wire n5923;
  wire [3:0] n5926;
  wire n5928;
  wire [15:0] n5929;
  reg [3:0] n5931;
  wire n5938;
  wire n5942;
  wire n5945;
  wire n5946;
  wire [1:0] n5947;
  wire [1:0] n5953;
  wire n5955;
  wire n5956;
  wire n5959;
  wire n5969;
  wire n5971;
  wire n5972;
  wire n5975;
  wire n5976;
  wire n5977;
  wire n5978;
  wire [3:0] n5979;
  wire [4:0] n5980;
  wire [4:0] n5981;
  wire [4:0] n5982;
  wire [4:0] n5983;
  wire n5985;
  wire [4:0] n5986;
  wire n5989;
  wire [31:0] n5990;
  wire n5992;
  wire [40:0] n5993;
  wire n5995;
  wire n5998;
  wire [3:0] n6000;
  wire n6001;
  reg n6002;
  wire n6003;
  reg n6004;
  wire [31:0] n6005;
  reg [31:0] n6006;
  wire [31:0] n6007;
  reg [31:0] n6008;
  wire [40:0] n6009;
  reg [40:0] n6010;
  wire n6012;
  wire n6013;
  wire n6014;
  wire [4:0] n6015;
  wire n6016;
  wire [30:0] n6017;
  wire [31:0] n6018;
  wire n6020;
  wire n6021;
  wire [30:0] n6022;
  wire [31:0] n6023;
  wire n6025;
  wire n6026;
  wire [39:0] n6027;
  wire [40:0] n6028;
  wire n6030;
  wire n6033;
  wire n6034;
  wire [3:0] n6035;
  wire n6036;
  reg n6037;
  wire n6038;
  reg n6039;
  wire [31:0] n6040;
  reg [31:0] n6041;
  wire [31:0] n6042;
  reg [31:0] n6043;
  wire [40:0] n6044;
  reg [40:0] n6045;
  wire n6047;
  wire [1:0] n6050;
  wire [1:0] n6051;
  wire [1:0] n6052;
  wire [64:0] n6053;
  wire n6054;
  wire n6055;
  wire n6056;
  wire n6057;
  wire n6058;
  wire n6059;
  wire n6060;
  wire n6061;
  wire [63:0] n6062;
  wire [63:0] n6063;
  wire [63:0] n6064;
  wire [40:0] n6065;
  wire [40:0] n6066;
  wire [66:0] n6067;
  wire [1:0] n6068;
  wire [63:0] n6069;
  wire [1:0] n6070;
  wire [1:0] n6071;
  wire n6072;
  wire n6073;
  wire n6074;
  wire [63:0] n6075;
  wire [63:0] n6076;
  wire [40:0] n6077;
  wire n6078;
  wire n6079;
  wire n6081;
  wire n6082;
  wire [4:0] n6083;
  wire n6084;
  wire n6086;
  wire n6087;
  wire n6089;
  wire n6090;
  wire n6092;
  wire n6093;
  wire [2:0] n6094;
  reg n6095;
  wire n6096;
  wire n6097;
  wire n6098;
  wire [71:0] n6100;
  wire [71:0] n6107;
  wire n6112;
  wire n6113;
  wire [1:0] n6116;
  wire [6:0] n6119;
  wire [31:0] n6120;
  wire [38:0] n6121;
  wire n6123;
  wire [1:0] n6129;
  wire [40:0] n6131;
  wire n6133;
  wire n6143;
  wire [4:0] n6144;
  wire n6146;
  wire n6147;
  wire n6148;
  wire n6149;
  wire n6150;
  wire n6151;
  wire [1:0] n6154;
  wire [1:0] n6155;
  wire [1:0] n6156;
  wire [1:0] n6157;
  wire [1:0] n6158;
  wire n6159;
  wire n6160;
  wire n6161;
  wire n6163;
  wire n6164;
  wire n6165;
  wire [4:0] n6166;
  wire n6168;
  wire n6169;
  wire n6171;
  wire n6172;
  wire n6173;
  wire n6175;
  wire n6176;
  wire n6177;
  wire n6178;
  wire n6179;
  wire n6180;
  wire [4:0] n6181;
  wire n6183;
  wire n6184;
  wire [6:0] n6185;
  wire [31:0] n6186;
  wire [1:0] n6187;
  wire n6189;
  wire [1:0] n6190;
  wire n6192;
  wire n6193;
  wire [1:0] n6194;
  wire [2:0] n6196;
  wire n6197;
  wire [2:0] n6198;
  wire [2:0] n6199;
  wire [38:0] n6200;
  wire n6201;
  wire [2:0] n6202;
  wire [2:0] n6203;
  wire [38:0] n6204;
  wire [38:0] n6205;
  wire [31:0] n6206;
  wire n6207;
  wire n6209;
  wire n6210;
  wire n6211;
  wire n6212;
  wire [1:0] n6213;
  wire [1:0] n6214;
  wire [31:0] n6215;
  wire [31:0] n6216;
  wire n6218;
  wire [76:0] n6219;
  wire [76:0] n6221;
  wire [1:0] n6224;
  wire [31:0] n6225;
  wire [6:0] n6226;
  reg [8:0] n6227;
  wire [13:0] n6228;
  wire [3:0] n6229;
  reg [3:0] n6230;
  reg [40:0] n6231;
  reg [71:0] n6232;
  wire [185:0] n6233;
  reg [1:0] n6234;
  wire [2:0] n6235;
  reg [76:0] n6236;
  reg n6237;
  wire [40:0] n6238;
  assign jtag_tdo_o = n6237; //(module output)
  assign \dmi_req_o_dmi_req_o[addr]  = n5767; //(module output)
  assign \dmi_req_o_dmi_req_o[op]  = n5768; //(module output)
  assign \dmi_req_o_dmi_req_o[data]  = n5769; //(module output)
  assign jtagspi_sck_o = n5809; //(module output)
  assign jtagspi_sdo_o = n5810; //(module output)
  assign jtagspi_csn_o = n5812; //(module output)
  assign n5767 = n6238[6:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:167:5  */
  assign n5768 = n6238[8:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:162:3  */
  assign n5769 = n6238[40:9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:81:3  */
  assign n5770 = {\dmi_rsp_i_dmi_rsp_i[ack] , \dmi_rsp_i_dmi_rsp_i[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:58:10  */
  assign tap_sync = n6228; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:63:10  */
  assign tap_ctrl_state = n6230; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:75:10  */
  assign tap_reg = n6233; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:82:10  */
  assign dr_trigger = n6235; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:94:10  */
  assign dmi_ctrl = n6236; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:102:16  */
  assign n5775 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:107:41  */
  assign n5780 = tap_sync[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:107:54  */
  assign n5781 = {n5780, jtag_tck_i};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:108:41  */
  assign n5782 = tap_sync[4:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:108:54  */
  assign n5783 = {n5782, jtag_tdi_i};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:109:41  */
  assign n5784 = tap_sync[7:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:109:54  */
  assign n5785 = {n5784, jtag_tms_i};
  assign n5786 = {n5785, n5783, n5781};
  assign n5789 = {3'b000, 3'b000, 3'b000};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:114:52  */
  assign n5793 = tap_sync[2:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:114:65  */
  assign n5795 = n5793 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:114:31  */
  assign n5796 = n5795 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:115:52  */
  assign n5799 = tap_sync[2:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:115:65  */
  assign n5801 = n5799 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:115:31  */
  assign n5802 = n5801 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:118:34  */
  assign n5804 = tap_sync[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:119:34  */
  assign n5805 = tap_sync[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:120:34  */
  assign n5806 = tap_sync[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:123:29  */
  assign n5807 = tap_sync[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:123:45  */
  assign n5808 = tap_reg[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:123:33  */
  assign n5809 = n5807 & n5808;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:124:29  */
  assign n5810 = tap_sync[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:125:32  */
  assign n5811 = tap_reg[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:125:20  */
  assign n5812 = ~n5811;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:131:16  */
  assign n5814 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:134:20  */
  assign n5816 = tap_sync[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:136:44  */
  assign n5817 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:136:48  */
  assign n5818 = ~n5817;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:136:31  */
  assign n5821 = n5818 ? 4'b1000 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:136:11  */
  assign n5823 = tap_ctrl_state == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:137:44  */
  assign n5824 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:137:48  */
  assign n5825 = ~n5824;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:137:31  */
  assign n5828 = n5825 ? 4'b1000 : 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:137:11  */
  assign n5830 = tap_ctrl_state == 4'b1000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:138:44  */
  assign n5831 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:138:48  */
  assign n5832 = ~n5831;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:138:31  */
  assign n5835 = n5832 ? 4'b0010 : 4'b1001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:138:11  */
  assign n5837 = tap_ctrl_state == 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:139:44  */
  assign n5838 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:139:48  */
  assign n5839 = ~n5838;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:139:31  */
  assign n5842 = n5839 ? 4'b0011 : 4'b0100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:139:11  */
  assign n5844 = tap_ctrl_state == 4'b0010;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:140:44  */
  assign n5845 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:140:48  */
  assign n5846 = ~n5845;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:140:31  */
  assign n5849 = n5846 ? 4'b0011 : 4'b0100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:140:11  */
  assign n5851 = tap_ctrl_state == 4'b0011;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:141:44  */
  assign n5852 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:141:48  */
  assign n5853 = ~n5852;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:141:31  */
  assign n5856 = n5853 ? 4'b0101 : 4'b0111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:141:11  */
  assign n5858 = tap_ctrl_state == 4'b0100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:142:44  */
  assign n5859 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:142:48  */
  assign n5860 = ~n5859;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:142:31  */
  assign n5863 = n5860 ? 4'b0101 : 4'b0110;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:142:11  */
  assign n5865 = tap_ctrl_state == 4'b0101;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:143:44  */
  assign n5866 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:143:48  */
  assign n5867 = ~n5866;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:143:31  */
  assign n5870 = n5867 ? 4'b0011 : 4'b0111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:143:11  */
  assign n5872 = tap_ctrl_state == 4'b0110;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:144:44  */
  assign n5873 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:144:48  */
  assign n5874 = ~n5873;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:144:31  */
  assign n5877 = n5874 ? 4'b1000 : 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:144:11  */
  assign n5879 = tap_ctrl_state == 4'b0111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:145:44  */
  assign n5880 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:145:48  */
  assign n5881 = ~n5880;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:145:31  */
  assign n5884 = n5881 ? 4'b1010 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:145:11  */
  assign n5886 = tap_ctrl_state == 4'b1001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:146:44  */
  assign n5887 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:146:48  */
  assign n5888 = ~n5887;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:146:31  */
  assign n5891 = n5888 ? 4'b1011 : 4'b1100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:146:11  */
  assign n5893 = tap_ctrl_state == 4'b1010;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:147:44  */
  assign n5894 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:147:48  */
  assign n5895 = ~n5894;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:147:31  */
  assign n5898 = n5895 ? 4'b1011 : 4'b1100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:147:11  */
  assign n5900 = tap_ctrl_state == 4'b1011;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:148:44  */
  assign n5901 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:148:48  */
  assign n5902 = ~n5901;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:148:31  */
  assign n5905 = n5902 ? 4'b1101 : 4'b1111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:148:11  */
  assign n5907 = tap_ctrl_state == 4'b1100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:149:44  */
  assign n5908 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:149:48  */
  assign n5909 = ~n5908;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:149:31  */
  assign n5912 = n5909 ? 4'b1101 : 4'b1110;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:149:11  */
  assign n5914 = tap_ctrl_state == 4'b1101;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:150:44  */
  assign n5915 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:150:48  */
  assign n5916 = ~n5915;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:150:31  */
  assign n5919 = n5916 ? 4'b1011 : 4'b1111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:150:11  */
  assign n5921 = tap_ctrl_state == 4'b1110;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:151:44  */
  assign n5922 = tap_sync[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:151:48  */
  assign n5923 = ~n5922;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:151:31  */
  assign n5926 = n5923 ? 4'b1000 : 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:151:11  */
  assign n5928 = tap_ctrl_state == 4'b1111;
  assign n5929 = {n5928, n5921, n5914, n5907, n5900, n5893, n5886, n5879, n5872, n5865, n5858, n5851, n5844, n5837, n5830, n5823};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:135:9  */
  always @*
    case (n5929)
      16'b1000000000000000: n5931 = n5926;
      16'b0100000000000000: n5931 = n5919;
      16'b0010000000000000: n5931 = n5912;
      16'b0001000000000000: n5931 = n5905;
      16'b0000100000000000: n5931 = n5898;
      16'b0000010000000000: n5931 = n5891;
      16'b0000001000000000: n5931 = n5884;
      16'b0000000100000000: n5931 = n5877;
      16'b0000000010000000: n5931 = n5870;
      16'b0000000001000000: n5931 = n5863;
      16'b0000000000100000: n5931 = n5856;
      16'b0000000000010000: n5931 = n5849;
      16'b0000000000001000: n5931 = n5842;
      16'b0000000000000100: n5931 = n5835;
      16'b0000000000000010: n5931 = n5828;
      16'b0000000000000001: n5931 = n5821;
      default: n5931 = 4'b0000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:161:16  */
  assign n5938 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:164:26  */
  assign n5942 = tap_ctrl_state == 4'b0111;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:164:7  */
  assign n5945 = n5942 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:169:44  */
  assign n5946 = dr_trigger[0]; // extract
  assign n5947 = {n5946, n5945};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:174:44  */
  assign n5953 = dr_trigger[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:174:49  */
  assign n5955 = n5953 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:174:27  */
  assign n5956 = n5955 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:181:16  */
  assign n5959 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:193:26  */
  assign n5969 = tap_ctrl_state == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:193:60  */
  assign n5971 = tap_ctrl_state == 4'b1010;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:193:41  */
  assign n5972 = n5969 | n5971;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:195:29  */
  assign n5975 = tap_ctrl_state == 4'b1011;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:195:55  */
  assign n5976 = tap_sync[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:195:41  */
  assign n5977 = n5976 & n5975;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:196:34  */
  assign n5978 = tap_sync[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:196:52  */
  assign n5979 = tap_reg[4:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:196:38  */
  assign n5980 = {n5978, n5979};
  assign n5981 = tap_reg[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:195:7  */
  assign n5982 = n5977 ? n5980 : n5981;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:193:7  */
  assign n5983 = n5972 ? 5'b00001 : n5982;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:200:26  */
  assign n5985 = tap_ctrl_state == 4'b0010;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:201:22  */
  assign n5986 = tap_reg[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:202:11  */
  assign n5989 = n5986 == 5'b00001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:203:59  */
  assign n5990 = tap_reg[103:72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:203:11  */
  assign n5992 = n5986 == 5'b10000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:204:59  */
  assign n5993 = tap_reg[185:145]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:204:11  */
  assign n5995 = n5986 == 5'b10001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:205:11  */
  assign n5998 = n5986 == 5'b10010;
  assign n6000 = {n5998, n5995, n5992, n5989};
  assign n6001 = tap_reg[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:201:9  */
  always @*
    case (n6000)
      4'b1000: n6002 = n6001;
      4'b0100: n6002 = n6001;
      4'b0010: n6002 = n6001;
      4'b0001: n6002 = n6001;
      default: n6002 = 1'b0;
    endcase
  assign n6003 = tap_reg[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:201:9  */
  always @*
    case (n6000)
      4'b1000: n6004 = 1'b1;
      4'b0100: n6004 = n6003;
      4'b0010: n6004 = n6003;
      4'b0001: n6004 = n6003;
      default: n6004 = n6003;
    endcase
  assign n6005 = tap_reg[39:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:201:9  */
  always @*
    case (n6000)
      4'b1000: n6006 = n6005;
      4'b0100: n6006 = n6005;
      4'b0010: n6006 = n6005;
      4'b0001: n6006 = 32'b00000000000000000000000000000001;
      default: n6006 = n6005;
    endcase
  assign n6007 = tap_reg[71:40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:201:9  */
  always @*
    case (n6000)
      4'b1000: n6008 = n6007;
      4'b0100: n6008 = n6007;
      4'b0010: n6008 = n5990;
      4'b0001: n6008 = n6007;
      default: n6008 = n6007;
    endcase
  assign n6009 = tap_reg[144:104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:201:9  */
  always @*
    case (n6000)
      4'b1000: n6010 = n6009;
      4'b0100: n6010 = n5993;
      4'b0010: n6010 = n6009;
      4'b0001: n6010 = n6009;
      default: n6010 = n6009;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:208:29  */
  assign n6012 = tap_ctrl_state == 4'b0011;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:208:55  */
  assign n6013 = tap_sync[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:208:41  */
  assign n6014 = n6013 & n6012;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:209:22  */
  assign n6015 = tap_reg[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:210:60  */
  assign n6016 = tap_sync[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:210:80  */
  assign n6017 = tap_reg[39:9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:210:64  */
  assign n6018 = {n6016, n6017};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:210:11  */
  assign n6020 = n6015 == 5'b00001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:211:60  */
  assign n6021 = tap_sync[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:211:79  */
  assign n6022 = tap_reg[71:41]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:211:64  */
  assign n6023 = {n6021, n6022};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:211:11  */
  assign n6025 = n6015 == 5'b10000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:212:60  */
  assign n6026 = tap_sync[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:212:77  */
  assign n6027 = tap_reg[144:105]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:212:64  */
  assign n6028 = {n6026, n6027};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:212:11  */
  assign n6030 = n6015 == 5'b10001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:213:11  */
  assign n6033 = n6015 == 5'b10010;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:214:60  */
  assign n6034 = tap_sync[12]; // extract
  assign n6035 = {n6033, n6030, n6025, n6020};
  assign n6036 = tap_reg[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:209:9  */
  always @*
    case (n6035)
      4'b1000: n6037 = n6036;
      4'b0100: n6037 = n6036;
      4'b0010: n6037 = n6036;
      4'b0001: n6037 = n6036;
      default: n6037 = n6034;
    endcase
  assign n6038 = tap_reg[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:209:9  */
  always @*
    case (n6035)
      4'b1000: n6039 = 1'b1;
      4'b0100: n6039 = n6038;
      4'b0010: n6039 = n6038;
      4'b0001: n6039 = n6038;
      default: n6039 = n6038;
    endcase
  assign n6040 = tap_reg[39:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:209:9  */
  always @*
    case (n6035)
      4'b1000: n6041 = n6040;
      4'b0100: n6041 = n6040;
      4'b0010: n6041 = n6040;
      4'b0001: n6041 = n6018;
      default: n6041 = n6040;
    endcase
  assign n6042 = tap_reg[71:40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:209:9  */
  always @*
    case (n6035)
      4'b1000: n6043 = n6042;
      4'b0100: n6043 = n6042;
      4'b0010: n6043 = n6023;
      4'b0001: n6043 = n6042;
      default: n6043 = n6042;
    endcase
  assign n6044 = tap_reg[144:104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:209:9  */
  always @*
    case (n6035)
      4'b1000: n6045 = n6044;
      4'b0100: n6045 = n6028;
      4'b0010: n6045 = n6044;
      4'b0001: n6045 = n6044;
      default: n6045 = n6044;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:216:29  */
  assign n6047 = tap_ctrl_state == 4'b0100;
  assign n6050 = {1'b0, 1'b0};
  assign n6051 = tap_reg[7:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:216:7  */
  assign n6052 = n6047 ? n6050 : n6051;
  assign n6053 = {n6043, n6041, n6039};
  assign n6054 = tap_reg[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:208:7  */
  assign n6055 = n6014 ? n6037 : n6054;
  assign n6056 = n6052[0]; // extract
  assign n6057 = tap_reg[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:208:7  */
  assign n6058 = n6014 ? n6057 : n6056;
  assign n6059 = n6052[1]; // extract
  assign n6060 = n6053[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:208:7  */
  assign n6061 = n6014 ? n6060 : n6059;
  assign n6062 = n6053[64:1]; // extract
  assign n6063 = tap_reg[71:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:208:7  */
  assign n6064 = n6014 ? n6062 : n6063;
  assign n6065 = tap_reg[144:104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:208:7  */
  assign n6066 = n6014 ? n6045 : n6065;
  assign n6067 = {n6064, n6061, n6058, n6055};
  assign n6068 = {n6004, n6002};
  assign n6069 = {n6008, n6006};
  assign n6070 = n6067[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:200:7  */
  assign n6071 = n5985 ? n6068 : n6070;
  assign n6072 = n6067[2]; // extract
  assign n6073 = tap_reg[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:200:7  */
  assign n6074 = n5985 ? n6073 : n6072;
  assign n6075 = n6067[66:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:200:7  */
  assign n6076 = n5985 ? n6069 : n6075;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:200:7  */
  assign n6077 = n5985 ? n6010 : n6066;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:222:19  */
  assign n6078 = tap_reg[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:224:23  */
  assign n6079 = tap_sync[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:225:28  */
  assign n6081 = tap_ctrl_state == 4'b1011;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:226:37  */
  assign n6082 = tap_reg[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:228:24  */
  assign n6083 = tap_reg[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:229:63  */
  assign n6084 = tap_reg[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:229:13  */
  assign n6086 = n6083 == 5'b00001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:230:62  */
  assign n6087 = tap_reg[40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:230:13  */
  assign n6089 = n6083 == 5'b10000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:231:60  */
  assign n6090 = tap_reg[104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:231:13  */
  assign n6092 = n6083 == 5'b10001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:232:57  */
  assign n6093 = tap_reg[5]; // extract
  assign n6094 = {n6092, n6089, n6086};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:228:11  */
  always @*
    case (n6094)
      3'b100: n6095 = n6090;
      3'b010: n6095 = n6087;
      3'b001: n6095 = n6084;
      default: n6095 = n6093;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:225:9  */
  assign n6096 = n6081 ? n6082 : n6095;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:224:7  */
  assign n6097 = n6079 ? n6096 : n6237;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:222:7  */
  assign n6098 = n6078 ? jtagspi_sdi_i : n6097;
  assign n6100 = {n6076, n6074, n6071, n5983};
  assign n6107 = {32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 1'b0, 1'b0, 1'b0, 5'b00000};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:242:47  */
  assign n6112 = dmi_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:243:47  */
  assign n6113 = dmi_ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:246:53  */
  assign n6116 = tap_reg[146:145]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:251:31  */
  assign n6119 = dmi_ctrl[76:70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:251:47  */
  assign n6120 = dmi_ctrl[37:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:251:36  */
  assign n6121 = {n6119, n6120};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:251:76  */
  assign n6123 = dmi_ctrl[5]; // extract
  assign n6129 = {n6123, n6123};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:251:53  */
  assign n6131 = {n6121, n6129};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:258:16  */
  assign n6133 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:269:22  */
  assign n6143 = dr_trigger[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:269:48  */
  assign n6144 = tap_reg[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:269:53  */
  assign n6146 = n6144 == 5'b10000;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:269:35  */
  assign n6147 = n6146 & n6143;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:270:47  */
  assign n6148 = tap_reg[56]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:271:47  */
  assign n6149 = tap_reg[57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:272:23  */
  assign n6150 = dmi_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:272:28  */
  assign n6151 = ~n6150;
  assign n6154 = {1'b0, 1'b0};
  assign n6155 = dmi_ctrl[4:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:272:7  */
  assign n6156 = n6151 ? n6154 : n6155;
  assign n6157 = {n6148, n6149};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:269:7  */
  assign n6158 = n6147 ? n6157 : n6156;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:278:20  */
  assign n6159 = dmi_ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:278:49  */
  assign n6160 = dmi_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:278:36  */
  assign n6161 = n6159 | n6160;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:280:23  */
  assign n6163 = dmi_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:280:51  */
  assign n6164 = dr_trigger[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:280:35  */
  assign n6165 = n6164 & n6163;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:280:77  */
  assign n6166 = tap_reg[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:280:82  */
  assign n6168 = n6166 == 5'b10001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:280:64  */
  assign n6169 = n6168 & n6165;
  assign n6171 = dmi_ctrl[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:280:7  */
  assign n6172 = n6169 ? 1'b1 : n6171;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:278:7  */
  assign n6173 = n6161 ? 1'b0 : n6172;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:286:20  */
  assign n6175 = dmi_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:286:25  */
  assign n6176 = ~n6175;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:287:22  */
  assign n6177 = dmi_ctrl[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:287:35  */
  assign n6178 = ~n6177;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:287:58  */
  assign n6179 = dr_trigger[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:287:42  */
  assign n6180 = n6179 & n6178;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:287:84  */
  assign n6181 = tap_reg[4:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:287:89  */
  assign n6183 = n6181 == 5'b10001;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:287:71  */
  assign n6184 = n6183 & n6180;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:288:40  */
  assign n6185 = tap_reg[144:138]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:289:40  */
  assign n6186 = tap_reg[137:106]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:290:26  */
  assign n6187 = tap_reg[105:104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:290:39  */
  assign n6189 = n6187 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:290:70  */
  assign n6190 = tap_reg[105:104]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:290:83  */
  assign n6192 = n6190 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:290:55  */
  assign n6193 = n6189 | n6192;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:291:41  */
  assign n6194 = tap_reg[105:104]; // extract
  assign n6196 = {n6194, 1'b1};
  assign n6197 = dmi_ctrl[0]; // extract
  assign n6198 = {2'b00, n6197};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:290:11  */
  assign n6199 = n6193 ? n6196 : n6198;
  assign n6200 = {n6185, n6186};
  assign n6201 = dmi_ctrl[0]; // extract
  assign n6202 = {2'b00, n6201};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:287:9  */
  assign n6203 = n6184 ? n6199 : n6202;
  assign n6204 = dmi_ctrl[76:38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:286:7  */
  assign n6205 = n6218 ? n6200 : n6204;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:296:37  */
  assign n6206 = n5770[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:297:23  */
  assign n6207 = n5770[32]; // extract
  assign n6209 = dmi_ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:297:9  */
  assign n6210 = n6207 ? 1'b0 : n6209;
  assign n6211 = n6203[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:286:7  */
  assign n6212 = n6176 ? n6211 : n6210;
  assign n6213 = n6203[2:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:286:7  */
  assign n6214 = n6176 ? n6213 : 2'b00;
  assign n6215 = dmi_ctrl[37:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:286:7  */
  assign n6216 = n6176 ? n6215 : n6206;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:286:7  */
  assign n6218 = n6184 & n6176;
  assign n6219 = {n6205, n6216, n6173, n6158, n6214, n6212};
  assign n6221 = {7'b0000000, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000, 1'b0, 1'b0, 1'b1, 2'b00, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:305:30  */
  assign n6224 = dmi_ctrl[2:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:306:30  */
  assign n6225 = dmi_ctrl[69:38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:307:30  */
  assign n6226 = dmi_ctrl[76:70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:106:5  */
  always @(posedge clk_i or posedge n5775)
    if (n5775)
      n6227 <= n5789;
    else
      n6227 <= n5786;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:102:5  */
  assign n6228 = {n5804, n5805, n5802, n5796, n5806, n6227};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:133:5  */
  assign n6229 = n5816 ? n5931 : tap_ctrl_state;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:133:5  */
  always @(posedge clk_i or posedge n5814)
    if (n5814)
      n6230 <= 4'b0000;
    else
      n6230 <= n6229;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:190:5  */
  always @(posedge clk_i or posedge n5959)
    if (n5959)
      n6231 <= 41'b00000000000000000000000000000000000000000;
    else
      n6231 <= n6077;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:190:5  */
  always @(posedge clk_i or posedge n5959)
    if (n5959)
      n6232 <= n6107;
    else
      n6232 <= n6100;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:181:5  */
  assign n6233 = {n6131, n6231, 14'b00000000000000, n6112, n6113, 1'b0, 3'b000, n6116, 6'b000111, 4'b0001, n6232};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:163:5  */
  always @(posedge clk_i or posedge n5938)
    if (n5938)
      n6234 <= 2'b00;
    else
      n6234 <= n5947;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:161:5  */
  assign n6235 = {n5956, n6234};
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:267:5  */
  always @(posedge clk_i or posedge n6133)
    if (n6133)
      n6236 <= n6221;
    else
      n6236 <= n6219;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:190:5  */
  always @(posedge clk_i or posedge n5959)
    if (n5959)
      n6237 <= 1'b0;
    else
      n6237 <= n6098;
  /* ../../ext/neorv32/rtl/core/neorv32_debug_dtm.vhd:181:5  */
  assign n6238 = {n6225, n6224, n6226};
endmodule

module neorv32_sysinfo_1_98304000_0_16384_16384_4_64_4_64_64_32_16_64_9e7924eaddd34398644d20f54977ca62b4d530f0
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] );
  wire [79:0] n5547;
  wire [31:0] n5549;
  wire n5550;
  wire n5551;
  wire [127:0] sysinfo;
  wire [1:0] buf_adr;
  wire buf_ack;
  wire n5553;
  wire n5556;
  wire n5557;
  wire n5558;
  wire [1:0] n5559;
  wire n5561;
  wire n5562;
  wire [31:0] n5563;
  wire n5578;
  wire n5582;
  wire n5586;
  wire n5590;
  wire n5594;
  wire n5598;
  wire n5602;
  wire n5607;
  wire n5611;
  wire n5615;
  wire n5619;
  wire n5623;
  wire n5627;
  wire n5631;
  wire n5635;
  wire n5639;
  wire n5643;
  wire n5647;
  wire n5651;
  wire n5655;
  wire n5659;
  wire n5663;
  wire n5667;
  wire n5671;
  wire n5675;
  wire n5679;
  wire n5684;
  wire n5688;
  wire n5692;
  wire n5696;
  wire [3:0] n5701;
  wire [3:0] n5706;
  wire [3:0] n5711;
  wire [3:0] n5716;
  wire [3:0] n5720;
  wire [3:0] n5724;
  wire [3:0] n5728;
  wire [3:0] n5732;
  wire n5735;
  wire n5737;
  wire n5738;
  wire [1:0] n5739;
  wire [1:0] n5750;
  wire [31:0] n5753;
  wire [31:0] n5756;
  wire [31:0] n5757;
  reg [31:0] n5758;
  wire [127:0] n5759;
  wire [1:0] n5760;
  reg [1:0] n5761;
  reg n5762;
  wire [33:0] n5763;
  wire [31:0] n5764;
  assign \bus_rsp_o_bus_rsp_o[data]  = n5549; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n5550; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n5551; //(module output)
  assign n5547 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n5549 = n5763[31:0]; // extract
  assign n5550 = n5763[32]; // extract
  assign n5551 = n5763[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:84:10  */
  assign sysinfo = n5759; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:87:10  */
  assign buf_adr = n5761; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:88:10  */
  assign buf_ack = n5762; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:97:16  */
  assign n5553 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:100:21  */
  assign n5556 = n5547[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:100:47  */
  assign n5557 = n5547[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:100:32  */
  assign n5558 = n5557 & n5556;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:100:76  */
  assign n5559 = n5547[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:100:89  */
  assign n5561 = n5559 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:100:57  */
  assign n5562 = n5561 & n5558;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:101:33  */
  assign n5563 = n5547[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:113:25  */
  assign n5578 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:114:25  */
  assign n5582 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:115:25  */
  assign n5586 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:116:25  */
  assign n5590 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:117:25  */
  assign n5594 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:118:25  */
  assign n5598 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:119:25  */
  assign n5602 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:121:25  */
  assign n5607 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:122:25  */
  assign n5611 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:123:25  */
  assign n5615 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:124:25  */
  assign n5619 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:125:25  */
  assign n5623 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:126:25  */
  assign n5627 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:127:25  */
  assign n5631 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:128:25  */
  assign n5635 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:129:25  */
  assign n5639 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:130:25  */
  assign n5643 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:131:25  */
  assign n5647 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:132:25  */
  assign n5651 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:133:25  */
  assign n5655 = 1'b1 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:134:25  */
  assign n5659 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:135:25  */
  assign n5663 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:136:25  */
  assign n5667 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:137:25  */
  assign n5671 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:138:25  */
  assign n5675 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:139:25  */
  assign n5679 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:141:25  */
  assign n5684 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:142:25  */
  assign n5688 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:143:25  */
  assign n5692 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:144:25  */
  assign n5696 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:147:98  */
  assign n5701 = 1'b0 ? 4'b0110 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:148:98  */
  assign n5706 = 1'b0 ? 4'b0010 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:150:98  */
  assign n5711 = 1'b0 ? 4'b0110 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:151:98  */
  assign n5716 = 1'b0 ? 4'b0010 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:153:101  */
  assign n5720 = 1'b1 ? 4'b0110 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:154:101  */
  assign n5724 = 1'b1 ? 4'b0100 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:156:102  */
  assign n5728 = 1'b0 ? 4'b0101 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:157:102  */
  assign n5732 = 1'b0 ? 4'b0110 : 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:164:16  */
  assign n5735 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:168:28  */
  assign n5737 = n5547[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:169:21  */
  assign n5738 = n5547[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:170:34  */
  assign n5739 = n5547[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:176:29  */
  assign n5750 = 2'b11 - buf_adr;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:176:60  */
  assign n5753 = buf_ack ? n5764 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:99:5  */
  assign n5756 = sysinfo[127:96]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:99:5  */
  assign n5757 = n5562 ? n5563 : n5756;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:99:5  */
  always @(posedge clk_i or posedge n5553)
    if (n5553)
      n5758 <= 32'b00000101110111000000000000000000;
    else
      n5758 <= n5757;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:97:5  */
  assign n5759 = {n5758, 8'b00000000, 8'b00000001, 8'b00001110, 8'b00001110, n5696, n5692, n5688, n5684, 1'b0, n5679, n5675, n5671, n5667, n5663, n5659, n5655, n5651, n5647, n5643, n5639, n5635, n5631, n5627, n5623, n5619, n5615, n5611, n5607, 1'b0, n5602, n5598, n5594, n5590, n5586, n5582, n5578, n5732, n5728, n5724, n5720, n5716, n5711, n5706, n5701};
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:167:5  */
  assign n5760 = n5738 ? n5739 : buf_adr;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:167:5  */
  always @(posedge clk_i or posedge n5735)
    if (n5735)
      n5761 <= 2'b00;
    else
      n5761 <= n5760;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:167:5  */
  always @(posedge clk_i or posedge n5735)
    if (n5735)
      n5762 <= 1'b0;
    else
      n5762 <= n5737;
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:164:5  */
  assign n5763 = {1'b0, buf_ack, n5753};
  /* ../../ext/neorv32/rtl/core/neorv32_sysinfo.vhd:176:29  */
  assign n5764 = sysinfo[n5750 * 32 +: 32]; //(Bmux)
endmodule

module neorv32_pwm_2
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   input  [7:0] clkgen_i,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output clkgen_en_o,
   output [15:0] pwm_o);
  wire [79:0] n5433;
  wire [31:0] n5435;
  wire n5436;
  wire n5437;
  wire [63:0] rdata;
  wire [31:0] rdata_sum;
  wire [1:0] sel;
  wire [1:0] we;
  wire [1:0] re;
  wire [1:0] ce;
  wire [1:0] pwm;
  wire n5441;
  wire n5443;
  wire [32:0] n5447;
  wire [32:0] n5448;
  wire [32:0] n5449;
  wire [33:0] n5451;
  wire [31:0] n5458;
  wire [31:0] n5460;
  wire [31:0] n5462;
  wire [31:0] n5463;
  wire n5465;
  wire n5466;
  wire [31:0] n5467;
  wire [31:0] pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5468;
  wire pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5469;
  wire pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5470;
  wire [3:0] n5478;
  wire n5480;
  wire n5481;
  wire n5483;
  wire n5484;
  wire n5485;
  wire n5486;
  wire n5487;
  wire n5488;
  wire n5489;
  wire n5490;
  wire n5491;
  wire n5492;
  wire n5493;
  wire n5494;
  wire n5495;
  wire [31:0] n5496;
  wire [31:0] pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5497;
  wire pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5498;
  wire pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5499;
  wire [3:0] n5507;
  wire n5509;
  wire n5510;
  wire n5512;
  wire n5513;
  wire n5514;
  wire n5515;
  wire n5516;
  wire n5517;
  wire n5518;
  wire n5519;
  wire n5520;
  wire n5521;
  wire n5522;
  localparam [15:0] n5524 = 16'b0000000000000000;
  wire [13:0] n5525;
  wire n5533;
  wire n5535;
  wire n5537;
  wire n5538;
  wire [63:0] n5539;
  wire [1:0] n5540;
  wire [1:0] n5541;
  wire [1:0] n5542;
  wire [1:0] n5543;
  wire [1:0] n5544;
  reg [33:0] n5545;
  wire [15:0] n5546;
  assign \bus_rsp_o_bus_rsp_o[data]  = n5435; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n5436; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n5437; //(module output)
  assign clkgen_en_o = n5538; //(module output)
  assign pwm_o = n5546; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:252:22  */
  assign n5433 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n5435 = n5545[31:0]; // extract
  assign n5436 = n5545[32]; // extract
  assign n5437 = n5545[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:56:10  */
  assign rdata = n5539; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:57:10  */
  assign rdata_sum = n5463; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:58:10  */
  assign sel = n5540; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:58:15  */
  assign we = n5541; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:58:19  */
  assign re = n5542; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:58:23  */
  assign ce = n5543; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:58:27  */
  assign pwm = n5544; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:66:16  */
  assign n5441 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:69:21  */
  assign n5443 = n5433[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:252:22  */
  assign n5447 = {1'b0, 32'b00000000000000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:241:3  */
  assign n5448 = {1'b1, rdata_sum};
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:69:7  */
  assign n5449 = n5443 ? n5448 : n5447;
  assign n5451 = {1'b0, n5449};
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:86:30  */
  assign n5458 = rdata[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:86:22  */
  assign n5460 = 32'b00000000000000000000000000000000 | n5458;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:86:30  */
  assign n5462 = rdata[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:86:22  */
  assign n5463 = n5460 | n5462;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:99:24  */
  assign n5465 = we[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:100:24  */
  assign n5466 = re[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:101:32  */
  assign n5467 = n5433[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:95:5  */
  neorv32_pwm_channel pwm_channel_gen_n1_neorv32_pwm_channel_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .we_i(n5465),
    .re_i(n5466),
    .wdata_i(n5467),
    .clkgen_i(clkgen_i),
    .rdata_o(pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5468),
    .clkgen_en_o(pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5469),
    .pwm_o(pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5470));
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:109:39  */
  assign n5478 = n5433[5:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:109:52  */
  assign n5480 = n5478 == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:109:19  */
  assign n5481 = n5480 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:18  */
  assign n5483 = sel[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:36  */
  assign n5484 = n5433[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:22  */
  assign n5485 = n5483 & n5484;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:59  */
  assign n5486 = n5433[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:40  */
  assign n5487 = n5485 & n5486;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:18  */
  assign n5488 = sel[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:36  */
  assign n5489 = n5433[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:22  */
  assign n5490 = n5488 & n5489;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:59  */
  assign n5491 = n5433[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:45  */
  assign n5492 = ~n5491;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:40  */
  assign n5493 = n5490 & n5492;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:99:24  */
  assign n5494 = we[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:100:24  */
  assign n5495 = re[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:101:32  */
  assign n5496 = n5433[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:95:5  */
  neorv32_pwm_channel pwm_channel_gen_n2_neorv32_pwm_channel_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .we_i(n5494),
    .re_i(n5495),
    .wdata_i(n5496),
    .clkgen_i(clkgen_i),
    .rdata_o(pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5497),
    .clkgen_en_o(pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5498),
    .pwm_o(pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5499));
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:109:39  */
  assign n5507 = n5433[5:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:109:52  */
  assign n5509 = n5507 == 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:109:19  */
  assign n5510 = n5509 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:18  */
  assign n5512 = sel[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:36  */
  assign n5513 = n5433[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:22  */
  assign n5514 = n5512 & n5513;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:59  */
  assign n5515 = n5433[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:110:40  */
  assign n5516 = n5514 & n5515;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:18  */
  assign n5517 = sel[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:36  */
  assign n5518 = n5433[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:22  */
  assign n5519 = n5517 & n5518;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:59  */
  assign n5520 = n5433[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:45  */
  assign n5521 = ~n5520;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:111:40  */
  assign n5522 = n5519 & n5521;
  assign n5525 = n5524[15:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n5533 = ce[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n5535 = 1'b0 | n5533;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n5537 = ce[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n5538 = n5535 | n5537;
  assign n5539 = {pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5468, pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5497};
  assign n5540 = {n5510, n5481};
  assign n5541 = {n5516, n5487};
  assign n5542 = {n5522, n5493};
  assign n5543 = {pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5498, pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5469};
  assign n5544 = {pwm_channel_gen_n2_neorv32_pwm_channel_inst_n5499, pwm_channel_gen_n1_neorv32_pwm_channel_inst_n5470};
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:68:5  */
  always @(posedge clk_i or posedge n5441)
    if (n5441)
      n5545 <= 34'b0000000000000000000000000000000000;
    else
      n5545 <= n5451;
  /* ../../ext/neorv32/rtl/core/neorv32_pwm.vhd:66:5  */
  assign n5546 = {n5525, pwm};
endmodule

module neorv32_twi_1
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   input  [7:0] clkgen_i,
   input  twi_sda_i,
   input  twi_scl_i,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output clkgen_en_o,
   output twi_sda_o,
   output twi_scl_o,
   output irq_o);
  wire [79:0] n5016;
  wire [31:0] n5018;
  wire n5019;
  wire n5020;
  wire [8:0] ctrl;
  wire [48:0] fifo;
  wire [17:0] clk_gen;
  wire [17:0] engine;
  wire [7:0] io_con;
  wire n5026;
  wire n5031;
  localparam [31:0] n5033 = 32'b00000000000000000000000000000000;
  wire n5034;
  wire n5035;
  wire n5036;
  wire n5037;
  wire n5038;
  wire [2:0] n5039;
  wire [3:0] n5040;
  wire n5041;
  wire [8:0] n5042;
  wire n5044;
  wire n5045;
  wire n5046;
  wire [2:0] n5047;
  wire [3:0] n5048;
  wire n5049;
  wire n5052;
  wire n5053;
  wire n5054;
  wire n5055;
  wire n5056;
  wire n5057;
  wire n5058;
  wire n5059;
  wire [8:0] n5060;
  wire [8:0] n5061;
  wire [4:0] n5062;
  wire [8:0] n5063;
  wire [3:0] n5064;
  wire [3:0] n5065;
  wire [4:0] n5066;
  wire [4:0] n5067;
  wire [8:0] n5068;
  wire [8:0] n5069;
  wire [3:0] n5070;
  wire [3:0] n5071;
  wire [4:0] n5072;
  wire [4:0] n5073;
  wire n5074;
  wire [8:0] n5075;
  wire [8:0] n5076;
  wire [3:0] n5077;
  wire [3:0] n5078;
  wire [4:0] n5079;
  wire [4:0] n5080;
  wire [5:0] n5083;
  wire [7:0] n5084;
  wire n5085;
  wire [33:0] n5086;
  wire [7:0] n5091;
  wire n5098;
  wire n5099;
  wire \tx_fifo_inst.half_o ;
  wire \tx_fifo_inst.free_o ;
  wire [10:0] \tx_fifo_inst.rdata_o ;
  wire \tx_fifo_inst.avail_o ;
  wire n5100;
  wire [10:0] n5101;
  wire n5102;
  wire n5104;
  wire n5108;
  wire n5109;
  wire n5110;
  wire n5111;
  wire n5112;
  wire n5113;
  wire [10:0] n5115;
  wire n5117;
  wire n5118;
  wire n5119;
  wire n5120;
  wire n5121;
  wire n5122;
  wire n5123;
  wire \rx_fifo_inst.half_o ;
  wire \rx_fifo_inst.free_o ;
  wire [8:0] \rx_fifo_inst.rdata_o ;
  wire \rx_fifo_inst.avail_o ;
  wire n5125;
  wire [8:0] n5126;
  wire n5127;
  wire n5129;
  wire n5132;
  wire [7:0] n5133;
  wire [8:0] n5134;
  wire n5135;
  wire n5137;
  wire n5138;
  wire n5139;
  wire n5140;
  wire n5141;
  wire n5142;
  wire n5143;
  wire n5146;
  wire n5148;
  wire n5149;
  wire n5150;
  wire n5151;
  wire n5152;
  wire n5153;
  wire n5154;
  wire n5160;
  wire n5164;
  wire n5165;
  wire [2:0] n5169;
  wire [3:0] n5173;
  wire [3:0] n5174;
  wire n5175;
  wire [3:0] n5178;
  wire [3:0] n5180;
  wire [4:0] n5181;
  wire [3:0] n5182;
  wire [3:0] n5183;
  wire n5184;
  wire n5185;
  wire [4:0] n5186;
  wire [3:0] n5187;
  wire [4:0] n5188;
  wire [4:0] n5189;
  wire [4:0] n5190;
  wire [4:0] n5191;
  wire [4:0] n5194;
  wire n5197;
  wire n5199;
  wire [3:0] n5203;
  wire n5204;
  wire n5205;
  wire n5206;
  wire n5207;
  wire n5208;
  wire n5210;
  wire n5211;
  wire n5212;
  wire n5213;
  wire [2:0] n5214;
  wire n5215;
  wire [3:0] n5216;
  wire [3:0] n5217;
  wire [3:0] n5218;
  wire [3:0] n5219;
  wire [7:0] n5220;
  wire [7:0] n5223;
  wire n5226;
  wire n5227;
  wire n5228;
  wire n5229;
  wire n5230;
  wire n5231;
  wire n5232;
  wire n5233;
  wire n5234;
  wire n5235;
  wire n5236;
  wire n5237;
  wire n5238;
  wire n5239;
  wire n5240;
  wire n5241;
  wire n5243;
  wire n5244;
  wire n5245;
  wire n5246;
  wire n5247;
  wire n5248;
  wire n5249;
  wire n5252;
  wire n5262;
  wire n5263;
  wire [1:0] n5264;
  wire n5265;
  wire n5266;
  wire [1:0] n5267;
  wire n5269;
  wire [2:0] n5270;
  wire [7:0] n5272;
  wire n5273;
  wire n5274;
  wire [8:0] n5275;
  wire n5276;
  wire n5277;
  wire n5278;
  wire [1:0] n5279;
  wire [1:0] n5280;
  wire [1:0] n5281;
  wire n5283;
  wire n5284;
  wire n5286;
  wire n5288;
  wire n5289;
  wire n5290;
  wire n5291;
  wire n5293;
  wire [1:0] n5296;
  wire [1:0] n5297;
  wire n5298;
  wire n5299;
  wire [1:0] n5300;
  wire [1:0] n5301;
  wire n5302;
  wire n5304;
  wire n5305;
  wire n5307;
  wire [1:0] n5310;
  wire [1:0] n5311;
  wire n5312;
  wire n5313;
  wire [1:0] n5314;
  wire [1:0] n5315;
  wire n5316;
  wire n5317;
  wire n5319;
  wire n5321;
  wire n5322;
  wire n5323;
  wire n5325;
  wire n5326;
  wire n5327;
  wire n5328;
  wire n5330;
  wire n5332;
  wire n5333;
  wire n5334;
  wire [3:0] n5335;
  wire n5337;
  wire n5338;
  wire n5339;
  wire n5341;
  wire n5342;
  wire n5343;
  wire n5344;
  wire n5345;
  wire n5346;
  wire [7:0] n5347;
  wire n5348;
  wire [8:0] n5349;
  wire [8:0] n5350;
  wire [8:0] n5351;
  wire n5352;
  wire [3:0] n5353;
  wire [3:0] n5355;
  wire [3:0] n5356;
  wire [3:0] n5357;
  wire [3:0] n5358;
  wire n5360;
  wire n5361;
  wire n5362;
  wire [1:0] n5365;
  wire [1:0] n5366;
  wire n5367;
  wire n5369;
  wire [3:0] n5373;
  reg [1:0] n5374;
  wire [3:0] n5375;
  reg [3:0] n5376;
  wire [8:0] n5377;
  reg [8:0] n5378;
  reg n5379;
  wire n5380;
  reg n5381;
  wire n5382;
  reg n5383;
  wire [16:0] n5384;
  wire [3:0] n5387;
  wire [1:0] n5388;
  wire [16:0] n5393;
  wire [3:0] n5395;
  wire [1:0] n5396;
  wire n5401;
  wire [1:0] n5402;
  wire n5404;
  wire n5405;
  wire n5406;
  wire n5408;
  wire n5409;
  wire n5410;
  wire n5411;
  wire n5412;
  wire n5413;
  wire n5414;
  reg n5415;
  wire [7:0] n5416;
  wire [7:0] n5417;
  wire [7:0] n5418;
  reg [7:0] n5419;
  wire [8:0] n5420;
  wire [48:0] n5421;
  reg [7:0] n5422;
  reg [4:0] n5423;
  wire [17:0] n5424;
  reg [16:0] n5425;
  wire [17:0] n5426;
  reg [1:0] n5427;
  reg [3:0] n5428;
  wire [7:0] n5429;
  reg [33:0] n5430;
  reg n5431;
  wire n5432;
  assign \bus_rsp_o_bus_rsp_o[data]  = n5018; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n5019; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n5020; //(module output)
  assign clkgen_en_o = n5197; //(module output)
  assign twi_sda_o = n5408; //(module output)
  assign twi_scl_o = n5409; //(module output)
  assign irq_o = n5431; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:366:23  */
  assign n5016 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:247:5  */
  assign n5018 = n5430[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:344:5  */
  assign n5019 = n5430[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:115:5  */
  assign n5020 = n5430[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:70:10  */
  assign ctrl = n5420; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:82:10  */
  assign fifo = n5421; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:93:10  */
  assign clk_gen = n5424; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:103:10  */
  assign engine = n5426; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:111:10  */
  assign io_con = n5429; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:119:16  */
  assign n5026 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:126:35  */
  assign n5031 = n5016[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:130:21  */
  assign n5034 = n5016[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:131:23  */
  assign n5035 = n5016[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:132:29  */
  assign n5036 = n5016[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:132:33  */
  assign n5037 = ~n5036;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:133:42  */
  assign n5038 = n5016[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:134:42  */
  assign n5039 = n5016[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:135:42  */
  assign n5040 = n5016[39:36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:136:42  */
  assign n5041 = n5016[40]; // extract
  assign n5042 = {n5041, n5040, n5039, n5038};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:139:29  */
  assign n5044 = n5016[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:139:33  */
  assign n5045 = ~n5044;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:140:70  */
  assign n5046 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:141:70  */
  assign n5047 = ctrl[3:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:142:70  */
  assign n5048 = ctrl[7:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:143:70  */
  assign n5049 = ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:147:65  */
  assign n5052 = io_con[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:148:65  */
  assign n5053 = io_con[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:149:58  */
  assign n5054 = fifo[48]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:149:49  */
  assign n5055 = ~n5054;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:150:54  */
  assign n5056 = fifo[45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:151:56  */
  assign n5057 = engine[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:151:69  */
  assign n5058 = fifo[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:151:61  */
  assign n5059 = n5057 | n5058;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:153:48  */
  assign n5060 = fifo[22:14]; // extract
  assign n5061 = {n5049, n5048, n5047, n5046};
  assign n5062 = {n5059, n5056, n5055, n5053, n5052};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:139:11  */
  assign n5063 = n5045 ? n5061 : n5060;
  assign n5064 = n5033[18:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:139:11  */
  assign n5065 = n5045 ? 4'b0000 : n5064;
  assign n5066 = n5033[31:27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:139:11  */
  assign n5067 = n5045 ? n5062 : n5066;
  assign n5068 = n5033[8:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:131:9  */
  assign n5069 = n5035 ? n5068 : n5063;
  assign n5070 = n5033[18:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:131:9  */
  assign n5071 = n5035 ? n5070 : n5065;
  assign n5072 = n5033[31:27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:131:9  */
  assign n5073 = n5035 ? n5072 : n5067;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:131:9  */
  assign n5074 = n5037 & n5035;
  assign n5075 = n5033[8:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:130:7  */
  assign n5076 = n5034 ? n5069 : n5075;
  assign n5077 = n5033[18:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:130:7  */
  assign n5078 = n5034 ? n5071 : n5077;
  assign n5079 = n5033[31:27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:130:7  */
  assign n5080 = n5034 ? n5073 : n5079;
  assign n5083 = n5033[14:9]; // extract
  assign n5084 = n5033[26:19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:130:7  */
  assign n5085 = n5074 & n5034;
  assign n5086 = {1'b0, n5031, n5080, n5084, n5078, n5083, n5076};
  assign n5091 = {4'b0000, 3'b000, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:165:26  */
  assign n5098 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:165:17  */
  assign n5099 = ~n5098;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:169:3  */
  neorv32_fifo_1_11_47ec8d98366433dc002e7721c9e37d5067547937 tx_fifo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n5100),
    .wdata_i(n5101),
    .we_i(n5102),
    .re_i(n5104),
    .half_o(),
    .free_o(\tx_fifo_inst.free_o ),
    .rdata_o(\tx_fifo_inst.rdata_o ),
    .avail_o(\tx_fifo_inst.avail_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:181:21  */
  assign n5100 = fifo[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:184:21  */
  assign n5101 = fifo[33:23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:185:21  */
  assign n5102 = fifo[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:188:21  */
  assign n5104 = fifo[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:193:40  */
  assign n5108 = n5016[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:193:66  */
  assign n5109 = n5016[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:193:51  */
  assign n5110 = n5109 & n5108;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:193:95  */
  assign n5111 = n5016[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:193:76  */
  assign n5112 = n5111 & n5110;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:193:24  */
  assign n5113 = n5112 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:194:34  */
  assign n5115 = n5016[42:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:195:37  */
  assign n5117 = engine[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:195:42  */
  assign n5118 = ~n5117;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:195:59  */
  assign n5119 = fifo[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:195:49  */
  assign n5120 = n5119 & n5118;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:195:88  */
  assign n5121 = clk_gen[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:195:75  */
  assign n5122 = n5121 & n5120;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:195:24  */
  assign n5123 = n5122 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:199:3  */
  neorv32_fifo_1_9_47ec8d98366433dc002e7721c9e37d5067547937 rx_fifo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n5125),
    .wdata_i(n5126),
    .we_i(n5127),
    .re_i(n5129),
    .half_o(),
    .free_o(\rx_fifo_inst.free_o ),
    .rdata_o(\rx_fifo_inst.rdata_o ),
    .avail_o(\rx_fifo_inst.avail_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:211:21  */
  assign n5125 = fifo[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:214:21  */
  assign n5126 = fifo[13:5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:215:21  */
  assign n5127 = fifo[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:218:21  */
  assign n5129 = fifo[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:223:31  */
  assign n5132 = engine[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:223:48  */
  assign n5133 = engine[15:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:223:35  */
  assign n5134 = {n5132, n5133};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:224:27  */
  assign n5135 = engine[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:225:40  */
  assign n5137 = n5016[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:225:66  */
  assign n5138 = n5016[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:225:69  */
  assign n5139 = ~n5138;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:225:51  */
  assign n5140 = n5139 & n5137;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:225:95  */
  assign n5141 = n5016[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:225:76  */
  assign n5142 = n5141 & n5140;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:225:24  */
  assign n5143 = n5142 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:231:16  */
  assign n5146 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:234:21  */
  assign n5148 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:234:42  */
  assign n5149 = fifo[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:234:33  */
  assign n5150 = ~n5149;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:234:28  */
  assign n5151 = n5148 & n5150;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:234:68  */
  assign n5152 = engine[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:234:57  */
  assign n5153 = ~n5152;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:234:52  */
  assign n5154 = n5151 & n5153;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:243:16  */
  assign n5160 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:247:16  */
  assign n5164 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:247:23  */
  assign n5165 = ~n5164;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:252:47  */
  assign n5169 = ctrl[3:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:253:23  */
  assign n5173 = clk_gen[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:253:34  */
  assign n5174 = ctrl[7:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:253:27  */
  assign n5175 = n5173 == n5174;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:257:63  */
  assign n5178 = clk_gen[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:257:68  */
  assign n5180 = n5178 + 4'b0001;
  assign n5181 = {1'b1, 4'b0000};
  assign n5182 = n5181[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:253:11  */
  assign n5183 = n5175 ? n5182 : n5180;
  assign n5184 = n5181[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:253:11  */
  assign n5185 = n5175 ? n5184 : 1'b0;
  assign n5186 = {n5185, n5183};
  assign n5187 = clk_gen[3:0]; // extract
  assign n5188 = {1'b0, n5187};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:252:9  */
  assign n5189 = n5432 ? n5186 : n5188;
  assign n5190 = {1'b0, 4'b0000};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:247:7  */
  assign n5191 = n5165 ? n5190 : n5189;
  assign n5194 = {1'b0, 4'b0000};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:265:23  */
  assign n5197 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:270:16  */
  assign n5199 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:274:39  */
  assign n5203 = clk_gen[9:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:275:16  */
  assign n5204 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:275:23  */
  assign n5205 = ~n5204;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:275:41  */
  assign n5206 = engine[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:275:46  */
  assign n5207 = ~n5206;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:275:30  */
  assign n5208 = n5205 | n5207;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:277:22  */
  assign n5210 = clk_gen[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:277:47  */
  assign n5211 = clk_gen[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:277:52  */
  assign n5212 = ~n5211;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:277:34  */
  assign n5213 = n5212 & n5210;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:278:47  */
  assign n5214 = clk_gen[8:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:278:79  */
  assign n5215 = clk_gen[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:278:60  */
  assign n5216 = {n5214, n5215};
  assign n5217 = clk_gen[9:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:277:7  */
  assign n5218 = n5213 ? n5216 : n5217;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:275:7  */
  assign n5219 = n5208 ? 4'b0001 : n5218;
  assign n5220 = {n5203, n5219};
  assign n5223 = {4'b0000, 4'b0000};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:284:43  */
  assign n5226 = clk_gen[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:284:73  */
  assign n5227 = clk_gen[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:284:52  */
  assign n5228 = ~n5227;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:284:47  */
  assign n5229 = n5226 & n5228;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:285:43  */
  assign n5230 = clk_gen[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:285:73  */
  assign n5231 = clk_gen[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:285:52  */
  assign n5232 = ~n5231;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:285:47  */
  assign n5233 = n5230 & n5232;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:286:43  */
  assign n5234 = clk_gen[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:286:73  */
  assign n5235 = clk_gen[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:286:52  */
  assign n5236 = ~n5235;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:286:47  */
  assign n5237 = n5234 & n5236;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:287:43  */
  assign n5238 = clk_gen[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:287:73  */
  assign n5239 = clk_gen[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:287:52  */
  assign n5240 = ~n5239;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:287:47  */
  assign n5241 = n5238 & n5240;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:291:36  */
  assign n5243 = io_con[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:291:72  */
  assign n5244 = io_con[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:291:76  */
  assign n5245 = ~n5244;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:291:51  */
  assign n5246 = n5245 & n5243;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:291:93  */
  assign n5247 = ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:291:83  */
  assign n5248 = n5247 & n5246;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:291:23  */
  assign n5249 = n5248 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:298:16  */
  assign n5252 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:309:43  */
  assign n5262 = io_con[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:309:56  */
  assign n5263 = io_con[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:309:47  */
  assign n5264 = {n5262, n5263};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:310:43  */
  assign n5265 = io_con[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:310:56  */
  assign n5266 = io_con[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:310:47  */
  assign n5267 = {n5265, n5266};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:316:31  */
  assign n5269 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:317:19  */
  assign n5270 = engine[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:322:41  */
  assign n5272 = fifo[41:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:322:92  */
  assign n5273 = fifo[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:322:75  */
  assign n5274 = ~n5273;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:322:72  */
  assign n5275 = {n5272, n5274};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:323:20  */
  assign n5276 = fifo[46]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:323:49  */
  assign n5277 = clk_gen[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:323:36  */
  assign n5278 = n5277 & n5276;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:324:54  */
  assign n5279 = fifo[44:43]; // extract
  assign n5280 = engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:323:11  */
  assign n5281 = n5278 ? n5279 : n5280;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:319:9  */
  assign n5283 = n5270 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:329:28  */
  assign n5284 = clk_gen[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:331:31  */
  assign n5286 = clk_gen[15]; // extract
  assign n5288 = io_con[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:331:11  */
  assign n5289 = n5286 ? 1'b0 : n5288;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:329:11  */
  assign n5290 = n5284 ? 1'b1 : n5289;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:335:28  */
  assign n5291 = clk_gen[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:337:31  */
  assign n5293 = clk_gen[17]; // extract
  assign n5296 = engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:337:11  */
  assign n5297 = n5293 ? 2'b00 : n5296;
  assign n5298 = io_con[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:337:11  */
  assign n5299 = n5293 ? 1'b0 : n5298;
  assign n5300 = engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:335:11  */
  assign n5301 = n5291 ? n5300 : n5297;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:335:11  */
  assign n5302 = n5291 ? 1'b1 : n5299;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:327:9  */
  assign n5304 = n5270 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:344:28  */
  assign n5305 = clk_gen[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:346:31  */
  assign n5307 = clk_gen[17]; // extract
  assign n5310 = engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:346:11  */
  assign n5311 = n5307 ? 2'b00 : n5310;
  assign n5312 = io_con[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:346:11  */
  assign n5313 = n5307 ? 1'b1 : n5312;
  assign n5314 = engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:344:11  */
  assign n5315 = n5305 ? n5314 : n5311;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:344:11  */
  assign n5316 = n5305 ? 1'b0 : n5313;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:351:28  */
  assign n5317 = clk_gen[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:353:31  */
  assign n5319 = clk_gen[15]; // extract
  assign n5321 = io_con[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:353:11  */
  assign n5322 = n5319 ? 1'b1 : n5321;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:351:11  */
  assign n5323 = n5317 ? 1'b0 : n5322;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:342:9  */
  assign n5325 = n5270 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:360:28  */
  assign n5326 = clk_gen[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:360:56  */
  assign n5327 = clk_gen[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:360:39  */
  assign n5328 = n5326 | n5327;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:362:31  */
  assign n5330 = clk_gen[15]; // extract
  assign n5332 = io_con[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:362:11  */
  assign n5333 = n5330 ? 1'b1 : n5332;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:360:11  */
  assign n5334 = n5328 ? 1'b0 : n5333;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:366:22  */
  assign n5335 = engine[6:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:366:29  */
  assign n5337 = n5335 == 4'b1001;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:366:57  */
  assign n5338 = clk_gen[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:366:39  */
  assign n5339 = n5338 & n5337;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:368:31  */
  assign n5341 = clk_gen[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:369:42  */
  assign n5342 = engine[15]; // extract
  assign n5343 = io_con[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:368:11  */
  assign n5344 = n5341 ? n5342 : n5343;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:366:11  */
  assign n5345 = n5339 ? 1'b0 : n5344;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:372:28  */
  assign n5346 = clk_gen[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:373:39  */
  assign n5347 = engine[14:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:373:70  */
  assign n5348 = io_con[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:373:52  */
  assign n5349 = {n5347, n5348};
  assign n5350 = engine[15:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:372:11  */
  assign n5351 = n5346 ? n5349 : n5350;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:376:28  */
  assign n5352 = clk_gen[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:377:64  */
  assign n5353 = engine[6:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:377:72  */
  assign n5355 = n5353 + 4'b0001;
  assign n5356 = engine[6:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:376:11  */
  assign n5357 = n5352 ? n5355 : n5356;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:380:22  */
  assign n5358 = engine[6:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:380:29  */
  assign n5360 = n5358 == 4'b1001;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:380:57  */
  assign n5361 = clk_gen[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:380:39  */
  assign n5362 = n5361 & n5360;
  assign n5365 = engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:380:11  */
  assign n5366 = n5362 ? 2'b00 : n5365;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:380:11  */
  assign n5367 = n5362 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:357:9  */
  assign n5369 = n5270 == 3'b111;
  assign n5373 = {n5369, n5325, n5304, n5283};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:317:7  */
  always @*
    case (n5373)
      4'b1000: n5374 = n5366;
      4'b0100: n5374 = n5315;
      4'b0010: n5374 = n5301;
      4'b0001: n5374 = n5281;
      default: n5374 = 2'b00;
    endcase
  assign n5375 = engine[6:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:317:7  */
  always @*
    case (n5373)
      4'b1000: n5376 = n5357;
      4'b0100: n5376 = n5375;
      4'b0010: n5376 = n5375;
      4'b0001: n5376 = 4'b0000;
      default: n5376 = n5375;
    endcase
  assign n5377 = engine[15:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:317:7  */
  always @*
    case (n5373)
      4'b1000: n5378 = n5351;
      4'b0100: n5378 = n5377;
      4'b0010: n5378 = n5377;
      4'b0001: n5378 = n5275;
      default: n5378 = n5377;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:317:7  */
  always @*
    case (n5373)
      4'b1000: n5379 = n5367;
      4'b0100: n5379 = 1'b0;
      4'b0010: n5379 = 1'b0;
      4'b0001: n5379 = 1'b0;
      default: n5379 = 1'b0;
    endcase
  assign n5380 = io_con[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:317:7  */
  always @*
    case (n5373)
      4'b1000: n5381 = n5345;
      4'b0100: n5381 = n5316;
      4'b0010: n5381 = n5290;
      4'b0001: n5381 = n5380;
      default: n5381 = 1'b1;
    endcase
  assign n5382 = io_con[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:317:7  */
  always @*
    case (n5373)
      4'b1000: n5383 = n5334;
      4'b0100: n5383 = n5323;
      4'b0010: n5383 = n5302;
      4'b0001: n5383 = n5382;
      default: n5383 = 1'b1;
    endcase
  assign n5384 = {n5379, n5378, n5376, n5269, n5374};
  assign n5387 = {n5267, n5264};
  assign n5388 = {n5383, n5381};
  assign n5393 = {1'b0, 9'b000000000, 4'b0000, 3'b000};
  assign n5395 = {2'b00, 2'b00};
  assign n5396 = {1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:396:40  */
  assign n5401 = engine[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:396:68  */
  assign n5402 = engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:396:81  */
  assign n5404 = n5402 != 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:396:51  */
  assign n5405 = n5404 & n5401;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:396:22  */
  assign n5406 = n5405 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:401:27  */
  assign n5408 = io_con[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:402:27  */
  assign n5409 = io_con[7]; // extract
  assign n5410 = n5042[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:117:3  */
  assign n5411 = ~n5026;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:117:3  */
  assign n5412 = n5085 & n5411;
  assign n5413 = ctrl[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:124:5  */
  assign n5414 = n5412 ? n5410 : n5413;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:124:5  */
  always @(posedge clk_i)
    n5415 <= n5414;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:119:5  */
  assign n5416 = n5042[7:0]; // extract
  assign n5417 = ctrl[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:124:5  */
  assign n5418 = n5085 ? n5416 : n5417;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:124:5  */
  always @(posedge clk_i or posedge n5026)
    if (n5026)
      n5419 <= n5091;
    else
      n5419 <= n5418;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:119:5  */
  assign n5420 = {n5415, n5419};
  assign n5421 = {\tx_fifo_inst.free_o , \rx_fifo_inst.free_o , \tx_fifo_inst.avail_o , \rx_fifo_inst.avail_o , \tx_fifo_inst.rdata_o , n5115, \rx_fifo_inst.rdata_o , n5134, n5123, n5143, n5113, n5135, n5099};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:273:5  */
  always @(posedge clk_i or posedge n5199)
    if (n5199)
      n5422 <= n5223;
    else
      n5422 <= n5220;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:246:5  */
  always @(posedge clk_i or posedge n5160)
    if (n5160)
      n5423 <= n5194;
    else
      n5423 <= n5191;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:243:5  */
  assign n5424 = {n5241, n5237, n5233, n5229, n5422, n5249, n5423};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:307:5  */
  always @(posedge clk_i or posedge n5252)
    if (n5252)
      n5425 <= n5393;
    else
      n5425 <= n5384;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:298:5  */
  assign n5426 = {n5406, n5425};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:307:5  */
  always @(posedge clk_i or posedge n5252)
    if (n5252)
      n5427 <= n5396;
    else
      n5427 <= n5388;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:307:5  */
  always @(posedge clk_i or posedge n5252)
    if (n5252)
      n5428 <= n5395;
    else
      n5428 <= n5387;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:298:5  */
  assign n5429 = {n5427, twi_scl_i, twi_sda_i, n5428};
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:124:5  */
  always @(posedge clk_i or posedge n5026)
    if (n5026)
      n5430 <= 34'b0000000000000000000000000000000000;
    else
      n5430 <= n5086;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:233:5  */
  always @(posedge clk_i or posedge n5146)
    if (n5146)
      n5431 <= 1'b0;
    else
      n5431 <= n5154;
  /* ../../ext/neorv32/rtl/core/neorv32_twi.vhd:252:22  */
  assign n5432 = clkgen_i[n5169 * 1 +: 1]; //(Bmux)
endmodule

module neorv32_spi_1
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   input  [7:0] clkgen_i,
   input  spi_dat_i,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output clkgen_en_o,
   output spi_clk_o,
   output spi_dat_o,
   output [7:0] spi_csn_o,
   output irq_o);
  wire [79:0] n4608;
  wire [31:0] n4610;
  wire n4611;
  wire n4612;
  wire [14:0] ctrl;
  wire [3:0] cdiv_cnt;
  wire spi_clk_en;
  wire [22:0] rtx_engine;
  wire [23:0] tx_fifo;
  wire [23:0] rx_fifo;
  wire n4619;
  wire n4631;
  localparam [31:0] n4633 = 32'b00000000000000000000000000000000;
  wire n4634;
  wire n4635;
  wire n4636;
  wire n4637;
  wire n4638;
  wire n4639;
  wire n4640;
  wire [2:0] n4641;
  wire [3:0] n4642;
  wire n4643;
  wire n4644;
  wire n4645;
  wire n4646;
  wire n4647;
  wire [14:0] n4648;
  wire n4650;
  wire n4651;
  wire n4652;
  wire n4653;
  wire n4654;
  wire [2:0] n4655;
  wire [3:0] n4656;
  wire n4657;
  wire n4658;
  wire n4659;
  wire n4660;
  wire n4661;
  wire n4662;
  wire n4663;
  wire n4664;
  wire n4665;
  wire n4666;
  wire n4667;
  wire n4668;
  wire n4671;
  wire n4672;
  wire n4673;
  wire n4674;
  wire [7:0] n4675;
  wire [10:0] n4676;
  wire [11:0] n4677;
  wire [1:0] n4678;
  wire [7:0] n4679;
  wire [7:0] n4680;
  wire [2:0] n4681;
  wire [2:0] n4682;
  wire [2:0] n4683;
  wire [11:0] n4684;
  wire [11:0] n4685;
  wire [1:0] n4686;
  wire [1:0] n4687;
  wire [10:0] n4688;
  wire [10:0] n4689;
  wire [10:0] n4690;
  wire [11:0] n4691;
  wire [11:0] n4692;
  wire [1:0] n4693;
  wire [1:0] n4694;
  wire n4695;
  wire [10:0] n4696;
  wire [10:0] n4697;
  wire [11:0] n4698;
  wire [11:0] n4699;
  wire [1:0] n4700;
  wire [1:0] n4701;
  wire [4:0] n4704;
  wire [1:0] n4705;
  wire n4706;
  wire [33:0] n4707;
  wire [14:0] n4712;
  wire \tx_fifo_inst.half_o ;
  wire \tx_fifo_inst.free_o ;
  wire [8:0] \tx_fifo_inst.rdata_o ;
  wire \tx_fifo_inst.avail_o ;
  wire n4715;
  wire [8:0] n4717;
  wire n4718;
  wire n4720;
  wire n4723;
  wire n4724;
  wire n4726;
  wire n4727;
  wire n4728;
  wire n4729;
  wire n4730;
  wire n4731;
  wire n4733;
  wire [7:0] n4734;
  wire [8:0] n4735;
  wire [2:0] n4737;
  wire n4739;
  wire n4740;
  wire \rx_fifo_inst.half_o ;
  wire \rx_fifo_inst.free_o ;
  wire [8:0] \rx_fifo_inst.rdata_o ;
  wire \rx_fifo_inst.avail_o ;
  wire n4742;
  wire [8:0] n4744;
  wire n4745;
  wire n4747;
  wire n4750;
  wire n4751;
  wire [7:0] n4752;
  wire [8:0] n4754;
  wire n4755;
  wire n4757;
  wire n4758;
  wire n4759;
  wire n4760;
  wire n4761;
  wire n4762;
  wire n4763;
  wire n4766;
  wire n4768;
  wire n4769;
  wire n4770;
  wire n4771;
  wire n4772;
  wire n4773;
  wire n4774;
  wire n4775;
  wire n4776;
  wire n4777;
  wire n4778;
  wire n4779;
  wire n4780;
  wire n4781;
  wire n4782;
  wire n4783;
  wire n4784;
  wire n4785;
  wire n4786;
  wire n4787;
  wire n4788;
  wire n4789;
  wire n4790;
  wire n4796;
  wire n4806;
  wire [2:0] n4807;
  wire n4808;
  wire n4810;
  wire n4811;
  wire [3:0] n4812;
  wire [7:0] n4813;
  wire [1:0] n4815;
  wire [1:0] n4816;
  wire [7:0] n4817;
  wire [7:0] n4818;
  wire [3:0] n4819;
  wire [3:0] n4820;
  wire [1:0] n4821;
  wire [1:0] n4822;
  wire [7:0] n4823;
  wire [7:0] n4824;
  wire n4826;
  wire n4828;
  wire n4829;
  wire n4830;
  wire n4831;
  wire n4832;
  wire n4833;
  wire [1:0] n4835;
  wire [1:0] n4836;
  wire n4838;
  wire n4840;
  wire n4841;
  wire n4842;
  wire n4843;
  wire n4844;
  wire [3:0] n4845;
  wire [3:0] n4847;
  wire [5:0] n4849;
  wire [1:0] n4850;
  wire [1:0] n4851;
  wire [5:0] n4852;
  wire [5:0] n4853;
  wire n4855;
  wire [6:0] n4856;
  wire n4857;
  wire [7:0] n4858;
  wire n4859;
  wire n4860;
  wire n4863;
  wire n4864;
  wire n4865;
  wire [1:0] n4867;
  wire n4868;
  wire n4869;
  wire [1:0] n4870;
  wire [1:0] n4871;
  wire [7:0] n4872;
  wire [7:0] n4873;
  wire n4874;
  wire n4875;
  wire n4876;
  wire n4878;
  wire n4879;
  wire [3:0] n4882;
  reg [1:0] n4883;
  wire [7:0] n4884;
  reg [7:0] n4885;
  wire [3:0] n4886;
  wire [3:0] n4887;
  reg [3:0] n4888;
  wire n4889;
  wire n4890;
  reg n4891;
  wire n4892;
  reg n4893;
  wire [3:0] n4894;
  reg [3:0] n4895;
  reg n4896;
  wire [2:0] n4897;
  wire [18:0] n4898;
  wire [18:0] n4903;
  wire [1:0] n4908;
  wire n4910;
  wire n4911;
  wire n4913;
  wire n4914;
  wire n4916;
  wire n4918;
  wire [2:0] n4919;
  localparam [7:0] n4922 = 8'b11111111;
  wire [7:0] n4926;
  wire n4933;
  wire n4935;
  wire n4936;
  wire [2:0] n4937;
  wire n4941;
  wire n4942;
  wire [3:0] n4943;
  wire n4944;
  wire [3:0] n4946;
  wire [3:0] n4948;
  wire n4951;
  wire [3:0] n4952;
  wire n4954;
  wire [3:0] n4956;
  wire n4958;
  wire n4967;
  wire [14:0] n4968;
  reg [14:0] n4969;
  reg [3:0] n4970;
  reg n4971;
  reg [18:0] n4972;
  reg [2:0] n4973;
  wire [22:0] n4974;
  wire [23:0] n4975;
  wire [23:0] n4976;
  reg [33:0] n4977;
  reg [7:0] n4978;
  reg n4979;
  wire n4980;
  wire n4981;
  wire n4982;
  wire n4983;
  wire n4984;
  wire n4985;
  wire n4986;
  wire n4987;
  wire n4988;
  wire n4989;
  wire n4990;
  wire n4991;
  wire n4992;
  wire n4993;
  wire n4994;
  wire n4995;
  wire n4996;
  wire n4997;
  wire n4998;
  wire n4999;
  wire n5000;
  wire n5001;
  wire n5002;
  wire n5003;
  wire n5004;
  wire n5005;
  wire n5006;
  wire n5007;
  wire n5008;
  wire n5009;
  wire n5010;
  wire n5011;
  wire n5012;
  wire n5013;
  wire [7:0] n5014;
  wire n5015;
  assign \bus_rsp_o_bus_rsp_o[data]  = n4610; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n4611; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n4612; //(module output)
  assign clkgen_en_o = n4967; //(module output)
  assign spi_clk_o = n4914; //(module output)
  assign spi_dat_o = n4913; //(module output)
  assign spi_csn_o = n4978; //(module output)
  assign irq_o = n4979; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:225:27  */
  assign n4608 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n4610 = n4977[31:0]; // extract
  assign n4611 = n4977[32]; // extract
  assign n4612 = n4977[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:81:10  */
  assign ctrl = n4969; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:84:10  */
  assign cdiv_cnt = n4970; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:85:10  */
  assign spi_clk_en = n4971; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:98:10  */
  assign rtx_engine = n4974; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:107:10  */
  assign tx_fifo = n4975; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:107:19  */
  assign rx_fifo = n4976; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:115:16  */
  assign n4619 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:129:35  */
  assign n4631 = n4608[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:134:21  */
  assign n4634 = n4608[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:135:23  */
  assign n4635 = n4608[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:136:29  */
  assign n4636 = n4608[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:136:33  */
  assign n4637 = ~n4636;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:137:48  */
  assign n4638 = n4608[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:138:48  */
  assign n4639 = n4608[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:139:48  */
  assign n4640 = n4608[34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:140:48  */
  assign n4641 = n4608[37:35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:141:48  */
  assign n4642 = n4608[41:38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:142:48  */
  assign n4643 = n4608[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:143:48  */
  assign n4644 = n4608[52]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:144:48  */
  assign n4645 = n4608[53]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:145:48  */
  assign n4646 = n4608[54]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:146:48  */
  assign n4647 = n4608[55]; // extract
  assign n4648 = {n4647, n4646, n4645, n4644, n4643, n4642, n4641, n4640, n4639, n4638};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:149:29  */
  assign n4650 = n4608[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:149:33  */
  assign n4651 = ~n4650;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:150:70  */
  assign n4652 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:151:70  */
  assign n4653 = ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:152:70  */
  assign n4654 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:153:70  */
  assign n4655 = ctrl[5:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:154:70  */
  assign n4656 = ctrl[9:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:155:70  */
  assign n4657 = ctrl[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:157:60  */
  assign n4658 = rx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:158:64  */
  assign n4659 = tx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:158:52  */
  assign n4660 = ~n4659;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:159:64  */
  assign n4661 = tx_fifo[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:159:52  */
  assign n4662 = ~n4661;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:160:64  */
  assign n4663 = tx_fifo[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:160:52  */
  assign n4664 = ~n4663;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:161:57  */
  assign n4665 = ctrl[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:162:57  */
  assign n4666 = ctrl[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:163:57  */
  assign n4667 = ctrl[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:164:57  */
  assign n4668 = ctrl[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:168:67  */
  assign n4671 = rtx_engine[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:169:60  */
  assign n4672 = rtx_engine[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:169:76  */
  assign n4673 = tx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:169:65  */
  assign n4674 = n4672 | n4673;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:171:56  */
  assign n4675 = rx_fifo[18:11]; // extract
  assign n4676 = {n4657, n4656, n4655, n4654, n4653, n4652};
  assign n4677 = {4'b0000, n4668, n4667, n4666, n4665, n4664, n4662, n4660, n4658};
  assign n4678 = {n4674, n4671};
  assign n4679 = n4676[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:149:11  */
  assign n4680 = n4651 ? n4679 : n4675;
  assign n4681 = n4676[10:8]; // extract
  assign n4682 = n4633[10:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:149:11  */
  assign n4683 = n4651 ? n4681 : n4682;
  assign n4684 = n4633[27:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:149:11  */
  assign n4685 = n4651 ? n4677 : n4684;
  assign n4686 = n4633[31:30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:149:11  */
  assign n4687 = n4651 ? n4678 : n4686;
  assign n4688 = {n4683, n4680};
  assign n4689 = n4633[10:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:135:9  */
  assign n4690 = n4635 ? n4689 : n4688;
  assign n4691 = n4633[27:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:135:9  */
  assign n4692 = n4635 ? n4691 : n4685;
  assign n4693 = n4633[31:30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:135:9  */
  assign n4694 = n4635 ? n4693 : n4687;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:135:9  */
  assign n4695 = n4637 & n4635;
  assign n4696 = n4633[10:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:134:7  */
  assign n4697 = n4634 ? n4690 : n4696;
  assign n4698 = n4633[27:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:134:7  */
  assign n4699 = n4634 ? n4692 : n4698;
  assign n4700 = n4633[31:30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:134:7  */
  assign n4701 = n4634 ? n4694 : n4700;
  assign n4704 = n4633[15:11]; // extract
  assign n4705 = n4633[29:28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:134:7  */
  assign n4706 = n4695 & n4634;
  assign n4707 = {1'b0, n4631, n4701, n4705, n4699, n4704, n4697};
  assign n4712 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 4'b0000, 3'b000, 1'b0, 1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:183:3  */
  neorv32_fifo_1_9_47ec8d98366433dc002e7721c9e37d5067547937 tx_fifo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n4715),
    .wdata_i(n4717),
    .we_i(n4718),
    .re_i(n4720),
    .half_o(\tx_fifo_inst.half_o ),
    .free_o(\tx_fifo_inst.free_o ),
    .rdata_o(\tx_fifo_inst.rdata_o ),
    .avail_o(\tx_fifo_inst.avail_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:195:24  */
  assign n4715 = tx_fifo[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:198:24  */
  assign n4717 = tx_fifo[10:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:199:24  */
  assign n4718 = tx_fifo[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:202:24  */
  assign n4720 = tx_fifo[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:207:29  */
  assign n4723 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:207:20  */
  assign n4724 = ~n4723;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:208:40  */
  assign n4726 = n4608[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:208:66  */
  assign n4727 = n4608[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:208:51  */
  assign n4728 = n4727 & n4726;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:208:95  */
  assign n4729 = n4608[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:208:76  */
  assign n4730 = n4729 & n4728;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:208:24  */
  assign n4731 = n4730 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:209:34  */
  assign n4733 = n4608[63]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:209:55  */
  assign n4734 = n4608[39:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:209:39  */
  assign n4735 = {n4733, n4734};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:210:41  */
  assign n4737 = rtx_engine[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:210:47  */
  assign n4739 = n4737 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:210:24  */
  assign n4740 = n4739 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:214:3  */
  neorv32_fifo_1_9_47ec8d98366433dc002e7721c9e37d5067547937 rx_fifo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n4742),
    .wdata_i(n4744),
    .we_i(n4745),
    .re_i(n4747),
    .half_o(\rx_fifo_inst.half_o ),
    .free_o(\rx_fifo_inst.free_o ),
    .rdata_o(\rx_fifo_inst.rdata_o ),
    .avail_o(\rx_fifo_inst.avail_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:226:24  */
  assign n4742 = rx_fifo[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:229:24  */
  assign n4744 = rx_fifo[10:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:230:24  */
  assign n4745 = rx_fifo[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:233:24  */
  assign n4747 = rx_fifo[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:238:29  */
  assign n4750 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:238:20  */
  assign n4751 = ~n4750;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:239:37  */
  assign n4752 = rtx_engine[11:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:239:24  */
  assign n4754 = {1'b0, n4752};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:240:31  */
  assign n4755 = rtx_engine[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:241:40  */
  assign n4757 = n4608[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:241:66  */
  assign n4758 = n4608[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:241:69  */
  assign n4759 = ~n4758;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:241:51  */
  assign n4760 = n4759 & n4757;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:241:95  */
  assign n4761 = n4608[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:241:76  */
  assign n4762 = n4761 & n4760;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:241:24  */
  assign n4763 = n4762 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:247:16  */
  assign n4766 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:250:21  */
  assign n4768 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:251:22  */
  assign n4769 = ctrl[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:251:52  */
  assign n4770 = rx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:251:35  */
  assign n4771 = n4769 & n4770;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:252:22  */
  assign n4772 = ctrl[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:252:52  */
  assign n4773 = tx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:252:40  */
  assign n4774 = ~n4773;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:252:35  */
  assign n4775 = n4772 & n4774;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:251:60  */
  assign n4776 = n4771 | n4775;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:253:22  */
  assign n4777 = ctrl[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:253:52  */
  assign n4778 = tx_fifo[23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:253:40  */
  assign n4779 = ~n4778;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:253:35  */
  assign n4780 = n4777 & n4779;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:252:60  */
  assign n4781 = n4776 | n4780;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:254:22  */
  assign n4782 = ctrl[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:254:52  */
  assign n4783 = tx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:254:40  */
  assign n4784 = ~n4783;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:254:35  */
  assign n4785 = n4782 & n4784;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:254:79  */
  assign n4786 = rtx_engine[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:254:64  */
  assign n4787 = ~n4786;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:254:59  */
  assign n4788 = n4785 & n4787;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:253:60  */
  assign n4789 = n4781 | n4788;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:250:28  */
  assign n4790 = n4768 & n4789;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:263:16  */
  assign n4796 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:276:35  */
  assign n4806 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:277:23  */
  assign n4807 = rtx_engine[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:281:37  */
  assign n4808 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:283:23  */
  assign n4810 = tx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:284:30  */
  assign n4811 = tx_fifo[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:285:50  */
  assign n4812 = tx_fifo[14:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:287:60  */
  assign n4813 = tx_fifo[18:11]; // extract
  assign n4815 = rtx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:284:13  */
  assign n4816 = n4811 ? n4815 : 2'b01;
  assign n4817 = rtx_engine[11:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:284:13  */
  assign n4818 = n4811 ? n4817 : n4813;
  assign n4819 = rtx_engine[21:18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:283:11  */
  assign n4820 = n4826 ? n4812 : n4819;
  assign n4821 = rtx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:283:11  */
  assign n4822 = n4810 ? n4816 : n4821;
  assign n4823 = rtx_engine[11:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:283:11  */
  assign n4824 = n4810 ? n4818 : n4823;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:283:11  */
  assign n4826 = n4811 & n4810;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:279:9  */
  assign n4828 = n4807 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:295:22  */
  assign n4829 = ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:296:42  */
  assign n4830 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:296:33  */
  assign n4831 = ~n4830;
  assign n4832 = rtx_engine[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:294:11  */
  assign n4833 = n4838 ? n4831 : n4832;
  assign n4835 = rtx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:294:11  */
  assign n4836 = spi_clk_en ? 2'b10 : n4835;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:294:11  */
  assign n4838 = n4829 & spi_clk_en;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:292:9  */
  assign n4840 = n4807 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:304:55  */
  assign n4841 = ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:304:69  */
  assign n4842 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:304:60  */
  assign n4843 = n4841 ^ n4842;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:304:45  */
  assign n4844 = ~n4843;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:306:83  */
  assign n4845 = rtx_engine[15:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:306:91  */
  assign n4847 = n4845 + 4'b0001;
  assign n4849 = {n4844, spi_dat_i, n4847};
  assign n4850 = rtx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:303:11  */
  assign n4851 = spi_clk_en ? 2'b11 : n4850;
  assign n4852 = rtx_engine[17:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:303:11  */
  assign n4853 = spi_clk_en ? n4849 : n4852;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:301:9  */
  assign n4855 = n4807 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:313:47  */
  assign n4856 = rtx_engine[10:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:313:73  */
  assign n4857 = rtx_engine[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:313:60  */
  assign n4858 = {n4856, n4857};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:314:34  */
  assign n4859 = rtx_engine[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:315:52  */
  assign n4860 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:319:52  */
  assign n4863 = ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:319:66  */
  assign n4864 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:319:57  */
  assign n4865 = n4863 ^ n4864;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:314:13  */
  assign n4867 = n4859 ? 2'b00 : 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:314:13  */
  assign n4868 = n4859 ? n4860 : n4865;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:312:11  */
  assign n4869 = n4876 ? 1'b1 : 1'b0;
  assign n4870 = rtx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:312:11  */
  assign n4871 = spi_clk_en ? n4867 : n4870;
  assign n4872 = rtx_engine[11:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:312:11  */
  assign n4873 = spi_clk_en ? n4858 : n4872;
  assign n4874 = rtx_engine[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:312:11  */
  assign n4875 = spi_clk_en ? n4868 : n4874;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:312:11  */
  assign n4876 = n4859 & spi_clk_en;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:310:9  */
  assign n4878 = n4807 == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:326:48  */
  assign n4879 = ctrl[2]; // extract
  assign n4882 = {n4878, n4855, n4840, n4828};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:277:7  */
  always @*
    case (n4882)
      4'b1000: n4883 = n4871;
      4'b0100: n4883 = n4851;
      4'b0010: n4883 = n4836;
      4'b0001: n4883 = n4822;
      default: n4883 = 2'b00;
    endcase
  assign n4884 = rtx_engine[11:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:277:7  */
  always @*
    case (n4882)
      4'b1000: n4885 = n4873;
      4'b0100: n4885 = n4884;
      4'b0010: n4885 = n4884;
      4'b0001: n4885 = n4824;
      default: n4885 = n4884;
    endcase
  assign n4886 = n4853[3:0]; // extract
  assign n4887 = rtx_engine[15:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:277:7  */
  always @*
    case (n4882)
      4'b1000: n4888 = n4887;
      4'b0100: n4888 = n4886;
      4'b0010: n4888 = n4887;
      4'b0001: n4888 = 4'b0000;
      default: n4888 = n4887;
    endcase
  assign n4889 = n4853[4]; // extract
  assign n4890 = rtx_engine[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:277:7  */
  always @*
    case (n4882)
      4'b1000: n4891 = n4890;
      4'b0100: n4891 = n4889;
      4'b0010: n4891 = n4890;
      4'b0001: n4891 = n4890;
      default: n4891 = n4890;
    endcase
  assign n4892 = n4853[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:277:7  */
  always @*
    case (n4882)
      4'b1000: n4893 = n4875;
      4'b0100: n4893 = n4892;
      4'b0010: n4893 = n4833;
      4'b0001: n4893 = n4808;
      default: n4893 = n4879;
    endcase
  assign n4894 = rtx_engine[21:18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:277:7  */
  always @*
    case (n4882)
      4'b1000: n4895 = n4894;
      4'b0100: n4895 = n4894;
      4'b0010: n4895 = n4894;
      4'b0001: n4895 = n4820;
      default: n4895 = 4'b0000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:277:7  */
  always @*
    case (n4882)
      4'b1000: n4896 = n4869;
      4'b0100: n4896 = 1'b0;
      4'b0010: n4896 = 1'b0;
      4'b0001: n4896 = 1'b0;
      default: n4896 = 1'b0;
    endcase
  assign n4897 = {n4806, n4883};
  assign n4898 = {n4896, n4895, n4893, n4891, n4888, n4885};
  assign n4903 = {1'b0, 4'b0000, 1'b0, 1'b0, 4'b0000, 8'b00000000};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:335:48  */
  assign n4908 = rtx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:335:61  */
  assign n4910 = n4908 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:335:26  */
  assign n4911 = n4910 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:338:31  */
  assign n4913 = rtx_engine[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:339:27  */
  assign n4914 = rtx_engine[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:344:16  */
  assign n4916 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:348:29  */
  assign n4918 = rtx_engine[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:57  */
  assign n4919 = rtx_engine[20:18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:348:7  */
  assign n4926 = n4918 ? n5014 : 8'b11111111;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:359:16  */
  assign n4933 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:364:16  */
  assign n4935 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:364:23  */
  assign n4936 = ~n4935;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:366:48  */
  assign n4937 = ctrl[5:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:366:72  */
  assign n4941 = ctrl[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:366:63  */
  assign n4942 = n5015 | n4941;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:367:29  */
  assign n4943 = ctrl[9:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:367:22  */
  assign n4944 = cdiv_cnt == n4943;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:371:60  */
  assign n4946 = cdiv_cnt + 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:367:9  */
  assign n4948 = n4944 ? 4'b0000 : n4946;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:367:9  */
  assign n4951 = n4944 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:366:7  */
  assign n4952 = n4942 ? n4948 : cdiv_cnt;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:366:7  */
  assign n4954 = n4942 ? n4951 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:364:7  */
  assign n4956 = n4936 ? 4'b0000 : n4952;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:364:7  */
  assign n4958 = n4936 ? 1'b0 : n4954;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:378:23  */
  assign n4967 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:127:5  */
  assign n4968 = n4706 ? n4648 : ctrl;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:127:5  */
  always @(posedge clk_i or posedge n4619)
    if (n4619)
      n4969 <= n4712;
    else
      n4969 <= n4968;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:362:5  */
  always @(posedge clk_i or posedge n4933)
    if (n4933)
      n4970 <= 4'b0000;
    else
      n4970 <= n4956;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:362:5  */
  always @(posedge clk_i or posedge n4933)
    if (n4933)
      n4971 <= 1'b0;
    else
      n4971 <= n4958;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:271:5  */
  always @(posedge clk_i or posedge n4796)
    if (n4796)
      n4972 <= n4903;
    else
      n4972 <= n4898;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:271:5  */
  always @(posedge clk_i or posedge n4796)
    if (n4796)
      n4973 <= 3'b000;
    else
      n4973 <= n4897;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:263:5  */
  assign n4974 = {n4972, n4911, n4973};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:263:5  */
  assign n4975 = {\tx_fifo_inst.half_o , n4724, \tx_fifo_inst.free_o , \tx_fifo_inst.avail_o , \tx_fifo_inst.rdata_o , n4735, n4740, n4731};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:359:5  */
  assign n4976 = {\rx_fifo_inst.half_o , n4751, \rx_fifo_inst.free_o , \rx_fifo_inst.avail_o , \rx_fifo_inst.rdata_o , n4754, n4763, n4755};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:127:5  */
  always @(posedge clk_i or posedge n4619)
    if (n4619)
      n4977 <= 34'b0000000000000000000000000000000000;
    else
      n4977 <= n4707;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:346:5  */
  always @(posedge clk_i or posedge n4916)
    if (n4916)
      n4978 <= 8'b11111111;
    else
      n4978 <= n4926;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:249:5  */
  always @(posedge clk_i or posedge n4766)
    if (n4766)
      n4979 <= 1'b0;
    else
      n4979 <= n4790;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4980 = n4919[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4981 = ~n4980;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4982 = n4919[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4983 = ~n4982;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4984 = n4981 & n4983;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4985 = n4981 & n4982;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4986 = n4980 & n4983;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4987 = n4980 & n4982;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4988 = n4919[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4989 = ~n4988;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4990 = n4984 & n4989;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4991 = n4984 & n4988;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4992 = n4985 & n4989;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4993 = n4985 & n4988;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4994 = n4986 & n4989;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4995 = n4986 & n4988;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4996 = n4987 & n4989;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4997 = n4987 & n4988;
  assign n4998 = n4922[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n4999 = n4990 ? 1'b0 : n4998;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:19  */
  assign n5000 = n4922[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n5001 = n4991 ? 1'b0 : n5000;
  assign n5002 = n4922[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n5003 = n4992 ? 1'b0 : n5002;
  assign n5004 = n4922[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n5005 = n4993 ? 1'b0 : n5004;
  assign n5006 = n4922[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n5007 = n4994 ? 1'b0 : n5006;
  assign n5008 = n4922[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n5009 = n4995 ? 1'b0 : n5008;
  assign n5010 = n4922[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n5011 = n4996 ? 1'b0 : n5010;
  assign n5012 = n4922[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:349:9  */
  assign n5013 = n4997 ? 1'b0 : n5012;
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:113:3  */
  assign n5014 = {n5013, n5011, n5009, n5007, n5005, n5003, n5001, n4999};
  /* ../../ext/neorv32/rtl/core/neorv32_spi.vhd:366:23  */
  assign n5015 = clkgen_i[n4937 * 1 +: 1]; //(Bmux)
endmodule

module neorv32_uart_1_1_e012e0243942cad1e54366b73ee6caff9501611d
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   input  [7:0] clkgen_i,
   input  uart_rxd_i,
   input  uart_cts_i,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output clkgen_en_o,
   output uart_txd_o,
   output uart_rts_o,
   output irq_rx_o,
   output irq_tx_o);
  wire [79:0] n4151;
  wire [31:0] n4153;
  wire n4154;
  wire n4155;
  wire uart_clk;
  wire [22:0] ctrl;
  wire [30:0] tx_engine;
  wire [29:0] rx_engine;
  wire [21:0] rx_fifo;
  wire [21:0] tx_fifo;
  wire n4162;
  wire n4176;
  localparam [31:0] n4178 = 32'b00000000000000000000000000000000;
  wire n4181;
  wire n4182;
  wire n4183;
  wire n4184;
  wire n4185;
  wire n4186;
  wire n4189;
  wire n4190;
  wire [2:0] n4191;
  wire [9:0] n4192;
  wire n4193;
  wire n4194;
  wire n4195;
  wire n4196;
  wire n4197;
  wire n4198;
  wire n4199;
  wire [22:0] n4200;
  wire [20:0] n4201;
  wire [22:0] n4202;
  wire [22:0] n4203;
  wire n4204;
  wire n4205;
  wire n4206;
  wire n4207;
  wire n4210;
  wire n4211;
  wire [2:0] n4212;
  wire [9:0] n4213;
  wire n4214;
  wire n4215;
  wire n4216;
  wire n4217;
  wire n4218;
  wire n4219;
  wire n4220;
  wire n4221;
  wire n4222;
  wire n4223;
  wire n4224;
  wire n4225;
  wire n4226;
  wire n4227;
  wire n4228;
  wire n4229;
  wire n4230;
  wire n4231;
  wire n4232;
  wire [7:0] n4233;
  wire [15:0] n4238;
  wire [26:0] n4239;
  wire [1:0] n4240;
  wire [15:0] n4241;
  wire [15:0] n4242;
  wire [10:0] n4243;
  wire [10:0] n4244;
  wire [10:0] n4245;
  wire [1:0] n4246;
  wire [1:0] n4247;
  wire [26:0] n4248;
  wire [26:0] n4249;
  wire [26:0] n4250;
  wire [1:0] n4251;
  wire [1:0] n4252;
  wire [20:0] n4253;
  wire [22:0] n4254;
  wire [22:0] n4255;
  wire [26:0] n4256;
  wire [26:0] n4257;
  wire [1:0] n4258;
  wire [1:0] n4259;
  wire [2:0] n4261;
  wire [20:0] n4262;
  wire [22:0] n4263;
  wire [22:0] n4264;
  wire [33:0] n4265;
  wire [22:0] n4270;
  wire n4273;
  wire [2:0] n4274;
  wire \tx_engine_fifo_inst.half_o ;
  wire \tx_engine_fifo_inst.free_o ;
  wire [7:0] \tx_engine_fifo_inst.rdata_o ;
  wire \tx_engine_fifo_inst.avail_o ;
  wire n4278;
  wire [7:0] n4280;
  wire n4281;
  wire n4283;
  wire n4287;
  wire n4288;
  wire n4289;
  wire n4290;
  wire n4291;
  wire n4292;
  wire n4293;
  wire [7:0] n4295;
  wire n4297;
  wire n4298;
  wire n4299;
  wire n4300;
  wire n4301;
  wire n4302;
  wire [2:0] n4305;
  wire n4307;
  wire n4308;
  wire n4311;
  wire n4313;
  wire n4314;
  wire n4315;
  wire n4316;
  wire n4317;
  wire n4318;
  wire n4319;
  wire n4320;
  wire n4321;
  wire n4322;
  wire n4323;
  wire \rx_engine_fifo_inst.half_o ;
  wire \rx_engine_fifo_inst.free_o ;
  wire [7:0] \rx_engine_fifo_inst.rdata_o ;
  wire \rx_engine_fifo_inst.avail_o ;
  wire n4328;
  wire [7:0] n4330;
  wire n4331;
  wire n4333;
  wire n4337;
  wire n4338;
  wire n4339;
  wire n4340;
  wire n4341;
  wire n4342;
  wire n4343;
  wire [7:0] n4345;
  wire n4346;
  wire n4348;
  wire n4349;
  wire n4350;
  wire n4351;
  wire n4352;
  wire n4353;
  wire n4354;
  wire n4357;
  wire n4359;
  wire n4360;
  wire n4361;
  wire n4362;
  wire n4363;
  wire n4364;
  wire n4365;
  wire n4366;
  wire n4367;
  wire n4368;
  wire n4369;
  wire n4370;
  wire n4371;
  wire n4372;
  wire n4378;
  wire n4387;
  wire [1:0] n4388;
  wire n4391;
  wire [2:0] n4392;
  wire [9:0] n4393;
  wire [7:0] n4395;
  wire [8:0] n4397;
  wire n4398;
  wire [1:0] n4400;
  wire [1:0] n4401;
  wire n4403;
  wire n4404;
  wire n4405;
  wire n4406;
  wire n4407;
  wire n4408;
  wire n4409;
  wire [1:0] n4411;
  wire [1:0] n4412;
  wire n4414;
  wire n4415;
  wire [9:0] n4416;
  wire n4418;
  wire [9:0] n4419;
  wire [3:0] n4420;
  wire [3:0] n4422;
  wire [7:0] n4423;
  wire [8:0] n4425;
  wire [9:0] n4426;
  wire [9:0] n4428;
  wire [22:0] n4429;
  wire [12:0] n4430;
  wire [12:0] n4431;
  wire [12:0] n4432;
  wire [9:0] n4433;
  wire [9:0] n4434;
  wire [22:0] n4435;
  wire [22:0] n4436;
  wire [22:0] n4437;
  wire [3:0] n4438;
  wire n4440;
  wire [1:0] n4443;
  wire [1:0] n4444;
  wire n4445;
  wire n4447;
  wire [2:0] n4449;
  reg [1:0] n4450;
  wire [8:0] n4451;
  wire [8:0] n4452;
  reg [8:0] n4453;
  wire [3:0] n4454;
  wire [3:0] n4455;
  reg [3:0] n4456;
  wire [9:0] n4457;
  wire [9:0] n4458;
  reg [9:0] n4459;
  reg n4460;
  reg n4461;
  wire [26:0] n4462;
  wire [2:0] n4463;
  wire [26:0] n4468;
  wire [2:0] n4469;
  wire [1:0] n4474;
  wire n4476;
  wire n4477;
  wire n4479;
  wire n4481;
  wire [1:0] n4489;
  wire [1:0] n4490;
  wire [1:0] n4491;
  wire n4493;
  wire [1:0] n4494;
  wire [8:0] n4495;
  wire [9:0] n4497;
  wire [1:0] n4499;
  wire n4501;
  wire n4503;
  wire n4504;
  wire n4506;
  wire [9:0] n4507;
  wire n4509;
  wire [9:0] n4510;
  wire [3:0] n4511;
  wire [3:0] n4513;
  wire n4514;
  wire [7:0] n4515;
  wire [8:0] n4516;
  wire [9:0] n4517;
  wire [9:0] n4519;
  wire [22:0] n4520;
  wire [12:0] n4521;
  wire [12:0] n4522;
  wire [12:0] n4523;
  wire [9:0] n4524;
  wire [9:0] n4525;
  wire [22:0] n4526;
  wire [22:0] n4527;
  wire [22:0] n4528;
  wire [3:0] n4529;
  wire n4531;
  wire n4534;
  wire n4535;
  wire n4536;
  wire n4538;
  wire [1:0] n4540;
  reg n4541;
  wire [8:0] n4542;
  wire [8:0] n4543;
  reg [8:0] n4544;
  wire [3:0] n4545;
  wire [3:0] n4546;
  reg [3:0] n4547;
  wire [9:0] n4548;
  wire [9:0] n4549;
  reg [9:0] n4550;
  reg n4551;
  wire [28:0] n4552;
  wire [28:0] n4555;
  wire n4559;
  wire n4562;
  wire n4563;
  wire n4565;
  wire n4566;
  wire n4567;
  wire n4568;
  wire n4570;
  wire n4571;
  wire n4572;
  wire n4578;
  wire n4580;
  wire n4581;
  wire n4582;
  wire n4583;
  wire n4584;
  wire n4587;
  wire n4589;
  reg [22:0] n4594;
  reg [2:0] n4595;
  reg [26:0] n4596;
  wire [30:0] n4597;
  reg n4598;
  reg [28:0] n4599;
  wire [29:0] n4600;
  wire [21:0] n4601;
  wire [21:0] n4602;
  reg [33:0] n4603;
  reg n4604;
  reg n4605;
  reg n4606;
  wire n4607;
  assign \bus_rsp_o_bus_rsp_o[data]  = n4153; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n4154; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n4155; //(module output)
  assign clkgen_en_o = n4273; //(module output)
  assign uart_txd_o = n4479; //(module output)
  assign uart_rts_o = n4604; //(module output)
  assign irq_rx_o = n4605; //(module output)
  assign irq_tx_o = n4606; //(module output)
  assign n4151 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n4153 = n4603[31:0]; // extract
  assign n4154 = n4603[32]; // extract
  assign n4155 = n4603[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:87:10  */
  assign uart_clk = n4607; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:104:10  */
  assign ctrl = n4594; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:117:10  */
  assign tx_engine = n4597; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:129:10  */
  assign rx_engine = n4600; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:142:10  */
  assign rx_fifo = n4601; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:142:19  */
  assign tx_fifo = n4602; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:150:16  */
  assign n4162 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:166:35  */
  assign n4176 = n4151[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:172:21  */
  assign n4181 = n4151[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:173:23  */
  assign n4182 = n4151[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:174:29  */
  assign n4183 = n4151[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:174:33  */
  assign n4184 = ~n4183;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:175:49  */
  assign n4185 = n4151[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:176:49  */
  assign n4186 = n4151[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:176:65  */
  assign n4189 = n4186 & 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:177:49  */
  assign n4190 = n4151[34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:178:49  */
  assign n4191 = n4151[37:35]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:179:49  */
  assign n4192 = n4151[47:38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:181:49  */
  assign n4193 = n4151[54]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:182:49  */
  assign n4194 = n4151[55]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:183:49  */
  assign n4195 = n4151[56]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:184:49  */
  assign n4196 = n4151[57]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:185:49  */
  assign n4197 = n4151[58]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:186:49  */
  assign n4198 = n4151[60]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:187:49  */
  assign n4199 = n4151[61]; // extract
  assign n4200 = {n4199, n4198, n4197, n4196, n4195, n4194, n4193, n4192, n4191, n4190, n4189, n4185};
  assign n4201 = ctrl[20:0]; // extract
  assign n4202 = {1'b0, 1'b0, n4201};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:174:11  */
  assign n4203 = n4184 ? n4200 : n4202;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:190:29  */
  assign n4204 = n4151[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:190:33  */
  assign n4205 = ~n4204;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:191:70  */
  assign n4206 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:192:70  */
  assign n4207 = ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:192:79  */
  assign n4210 = n4207 & 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:193:70  */
  assign n4211 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:194:70  */
  assign n4212 = ctrl[5:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:195:70  */
  assign n4213 = ctrl[15:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:197:73  */
  assign n4214 = rx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:198:73  */
  assign n4215 = rx_fifo[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:199:77  */
  assign n4216 = rx_fifo[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:199:65  */
  assign n4217 = ~n4216;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:200:77  */
  assign n4218 = tx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:200:65  */
  assign n4219 = ~n4218;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:201:77  */
  assign n4220 = tx_fifo[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:201:65  */
  assign n4221 = ~n4220;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:202:77  */
  assign n4222 = tx_fifo[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:202:65  */
  assign n4223 = ~n4222;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:204:70  */
  assign n4224 = ctrl[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:205:70  */
  assign n4225 = ctrl[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:206:70  */
  assign n4226 = ctrl[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:207:70  */
  assign n4227 = ctrl[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:208:70  */
  assign n4228 = ctrl[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:210:75  */
  assign n4229 = rx_engine[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:211:75  */
  assign n4230 = tx_engine[27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:211:91  */
  assign n4231 = tx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:211:80  */
  assign n4232 = n4230 | n4231;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:213:91  */
  assign n4233 = rx_fifo[18:11]; // extract
  assign n4238 = {4'b0000, 4'b0000, n4233};
  assign n4239 = {n4228, n4227, n4226, n4225, n4224, n4223, n4221, n4219, n4217, n4215, n4214, n4213, n4212, n4211, n4210, n4206};
  assign n4240 = {n4232, n4229};
  assign n4241 = n4239[15:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:190:11  */
  assign n4242 = n4205 ? n4241 : n4238;
  assign n4243 = n4239[26:16]; // extract
  assign n4244 = n4178[26:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:190:11  */
  assign n4245 = n4205 ? n4243 : n4244;
  assign n4246 = n4178[31:30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:190:11  */
  assign n4247 = n4205 ? n4240 : n4246;
  assign n4248 = {n4245, n4242};
  assign n4249 = n4178[26:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:173:9  */
  assign n4250 = n4182 ? n4249 : n4248;
  assign n4251 = n4178[31:30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:173:9  */
  assign n4252 = n4182 ? n4251 : n4247;
  assign n4253 = ctrl[20:0]; // extract
  assign n4254 = {1'b0, 1'b0, n4253};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:173:9  */
  assign n4255 = n4182 ? n4203 : n4254;
  assign n4256 = n4178[26:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:172:7  */
  assign n4257 = n4181 ? n4250 : n4256;
  assign n4258 = n4178[31:30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:172:7  */
  assign n4259 = n4181 ? n4252 : n4258;
  assign n4261 = n4178[29:27]; // extract
  assign n4262 = ctrl[20:0]; // extract
  assign n4263 = {1'b0, 1'b0, n4262};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:172:7  */
  assign n4264 = n4181 ? n4255 : n4263;
  assign n4265 = {1'b0, n4176, n4259, n4261, n4257};
  assign n4270 = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 10'b0000000000, 3'b000, 1'b0, 1'b0, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:224:23  */
  assign n4273 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:225:52  */
  assign n4274 = ctrl[5:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:230:3  */
  neorv32_fifo_1_8_47ec8d98366433dc002e7721c9e37d5067547937 tx_engine_fifo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n4278),
    .wdata_i(n4280),
    .we_i(n4281),
    .re_i(n4283),
    .half_o(\tx_engine_fifo_inst.half_o ),
    .free_o(\tx_engine_fifo_inst.free_o ),
    .rdata_o(\tx_engine_fifo_inst.rdata_o ),
    .avail_o(\tx_engine_fifo_inst.avail_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:242:24  */
  assign n4278 = tx_fifo[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:244:24  */
  assign n4280 = tx_fifo[10:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:245:24  */
  assign n4281 = tx_fifo[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:247:24  */
  assign n4283 = tx_fifo[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:252:35  */
  assign n4287 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:252:42  */
  assign n4288 = ~n4287;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:252:58  */
  assign n4289 = ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:252:49  */
  assign n4290 = n4288 | n4289;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:252:83  */
  assign n4291 = ctrl[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:252:74  */
  assign n4292 = n4290 | n4291;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:252:24  */
  assign n4293 = n4292 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:253:34  */
  assign n4295 = n4151[39:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:254:40  */
  assign n4297 = n4151[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:254:66  */
  assign n4298 = n4151[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:254:51  */
  assign n4299 = n4298 & n4297;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:254:95  */
  assign n4300 = n4151[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:254:76  */
  assign n4301 = n4300 & n4299;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:254:24  */
  assign n4302 = n4301 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:255:40  */
  assign n4305 = tx_engine[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:255:46  */
  assign n4307 = n4305 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:255:24  */
  assign n4308 = n4307 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:260:16  */
  assign n4311 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:263:24  */
  assign n4313 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:264:25  */
  assign n4314 = ctrl[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:264:55  */
  assign n4315 = tx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:264:43  */
  assign n4316 = ~n4315;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:264:38  */
  assign n4317 = n4314 & n4316;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:265:25  */
  assign n4318 = ctrl[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:265:55  */
  assign n4319 = tx_fifo[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:265:43  */
  assign n4320 = ~n4319;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:265:38  */
  assign n4321 = n4318 & n4320;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:264:63  */
  assign n4322 = n4317 | n4321;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:263:31  */
  assign n4323 = n4313 & n4322;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:272:3  */
  neorv32_fifo_1_8_47ec8d98366433dc002e7721c9e37d5067547937 rx_engine_fifo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .clear_i(n4328),
    .wdata_i(n4330),
    .we_i(n4331),
    .re_i(n4333),
    .half_o(\rx_engine_fifo_inst.half_o ),
    .free_o(\rx_engine_fifo_inst.free_o ),
    .rdata_o(\rx_engine_fifo_inst.rdata_o ),
    .avail_o(\rx_engine_fifo_inst.avail_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:283:24  */
  assign n4328 = rx_fifo[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:285:24  */
  assign n4330 = rx_fifo[10:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:286:24  */
  assign n4331 = rx_fifo[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:288:24  */
  assign n4333 = rx_fifo[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:293:35  */
  assign n4337 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:293:42  */
  assign n4338 = ~n4337;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:293:58  */
  assign n4339 = ctrl[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:293:49  */
  assign n4340 = n4338 | n4339;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:293:83  */
  assign n4341 = ctrl[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:293:74  */
  assign n4342 = n4340 | n4341;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:293:24  */
  assign n4343 = n4342 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:294:34  */
  assign n4345 = rx_engine[9:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:295:30  */
  assign n4346 = rx_engine[25]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:296:40  */
  assign n4348 = n4151[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:296:66  */
  assign n4349 = n4151[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:296:69  */
  assign n4350 = ~n4349;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:296:51  */
  assign n4351 = n4350 & n4348;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:296:95  */
  assign n4352 = n4151[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:296:76  */
  assign n4353 = n4352 & n4351;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:296:24  */
  assign n4354 = n4353 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:301:16  */
  assign n4357 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:304:24  */
  assign n4359 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:305:25  */
  assign n4360 = ctrl[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:305:51  */
  assign n4361 = rx_fifo[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:305:39  */
  assign n4362 = n4360 & n4361;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:306:25  */
  assign n4363 = ctrl[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:306:51  */
  assign n4364 = rx_fifo[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:306:39  */
  assign n4365 = n4363 & n4364;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:305:58  */
  assign n4366 = n4362 | n4365;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:307:25  */
  assign n4367 = ctrl[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:307:56  */
  assign n4368 = rx_fifo[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:307:44  */
  assign n4369 = ~n4368;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:307:39  */
  assign n4370 = n4367 & n4369;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:306:58  */
  assign n4371 = n4366 | n4370;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:304:31  */
  assign n4372 = n4359 & n4371;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:316:16  */
  assign n4378 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:326:47  */
  assign n4387 = tx_engine[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:326:51  */
  assign n4388 = {n4387, uart_cts_i};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:333:34  */
  assign n4391 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:334:22  */
  assign n4392 = tx_engine[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:338:37  */
  assign n4393 = ctrl[15:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:340:40  */
  assign n4395 = tx_fifo[18:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:340:46  */
  assign n4397 = {n4395, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:341:23  */
  assign n4398 = tx_fifo[20]; // extract
  assign n4400 = tx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:341:11  */
  assign n4401 = n4398 ? 2'b01 : n4400;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:336:9  */
  assign n4403 = n4392 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:348:34  */
  assign n4404 = tx_engine[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:348:38  */
  assign n4405 = ~n4404;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:348:54  */
  assign n4406 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:348:62  */
  assign n4407 = ~n4406;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:348:45  */
  assign n4408 = n4405 | n4407;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:347:31  */
  assign n4409 = n4408 & uart_clk;
  assign n4411 = tx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:347:11  */
  assign n4412 = n4409 ? 2'b11 : n4411;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:345:9  */
  assign n4414 = n4392 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:354:42  */
  assign n4415 = tx_engine[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:356:27  */
  assign n4416 = tx_engine[25:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:356:35  */
  assign n4418 = n4416 == 10'b0000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:357:41  */
  assign n4419 = ctrl[15:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:358:73  */
  assign n4420 = tx_engine[15:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:358:81  */
  assign n4422 = n4420 - 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:359:56  */
  assign n4423 = tx_engine[11:4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:359:40  */
  assign n4425 = {1'b1, n4423};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:361:73  */
  assign n4426 = tx_engine[25:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:361:82  */
  assign n4428 = n4426 - 10'b0000000001;
  assign n4429 = {n4419, n4422, n4425};
  assign n4430 = n4429[12:0]; // extract
  assign n4431 = tx_engine[15:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:356:13  */
  assign n4432 = n4418 ? n4430 : n4431;
  assign n4433 = n4429[22:13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:356:13  */
  assign n4434 = n4418 ? n4433 : n4428;
  assign n4435 = {n4434, n4432};
  assign n4436 = tx_engine[25:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:355:11  */
  assign n4437 = uart_clk ? n4435 : n4436;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:364:25  */
  assign n4438 = tx_engine[15:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:364:32  */
  assign n4440 = n4438 == 4'b0000;
  assign n4443 = tx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:364:11  */
  assign n4444 = n4440 ? 2'b00 : n4443;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:364:11  */
  assign n4445 = n4440 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:352:9  */
  assign n4447 = n4392 == 3'b111;
  assign n4449 = {n4447, n4414, n4403};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:334:7  */
  always @*
    case (n4449)
      3'b100: n4450 = n4444;
      3'b010: n4450 = n4412;
      3'b001: n4450 = n4401;
      default: n4450 = 2'b00;
    endcase
  assign n4451 = n4437[8:0]; // extract
  assign n4452 = tx_engine[11:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:334:7  */
  always @*
    case (n4449)
      3'b100: n4453 = n4451;
      3'b010: n4453 = n4452;
      3'b001: n4453 = n4397;
      default: n4453 = n4452;
    endcase
  assign n4454 = n4437[12:9]; // extract
  assign n4455 = tx_engine[15:12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:334:7  */
  always @*
    case (n4449)
      3'b100: n4456 = n4454;
      3'b010: n4456 = n4455;
      3'b001: n4456 = 4'b1011;
      default: n4456 = n4455;
    endcase
  assign n4457 = n4437[22:13]; // extract
  assign n4458 = tx_engine[25:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:334:7  */
  always @*
    case (n4449)
      3'b100: n4459 = n4457;
      3'b010: n4459 = n4458;
      3'b001: n4459 = n4393;
      default: n4459 = n4458;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:334:7  */
  always @*
    case (n4449)
      3'b100: n4460 = n4445;
      3'b010: n4460 = 1'b0;
      3'b001: n4460 = 1'b0;
      default: n4460 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:334:7  */
  always @*
    case (n4449)
      3'b100: n4461 = n4415;
      3'b010: n4461 = 1'b1;
      3'b001: n4461 = 1'b1;
      default: n4461 = 1'b1;
    endcase
  assign n4462 = {n4460, n4459, n4456, n4453, n4391, n4450};
  assign n4463 = {n4461, n4388};
  assign n4468 = {1'b0, 10'b0000000000, 4'b0000, 9'b000000000, 3'b000};
  assign n4469 = {1'b1, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:378:46  */
  assign n4474 = tx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:378:59  */
  assign n4476 = n4474 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:378:25  */
  assign n4477 = n4476 ? 1'b0 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:381:27  */
  assign n4479 = tx_engine[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:388:16  */
  assign n4481 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:399:53  */
  assign n4489 = rx_engine[28:27]; // extract
  assign n4490 = rx_engine[27:26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:398:7  */
  assign n4491 = uart_clk ? n4489 : n4490;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:406:34  */
  assign n4493 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:407:22  */
  assign n4494 = rx_engine[1:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:411:47  */
  assign n4495 = ctrl[15:7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:411:36  */
  assign n4497 = {1'b0, n4495};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:413:29  */
  assign n4499 = rx_engine[27:26]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:413:42  */
  assign n4501 = n4499 == 2'b01;
  assign n4503 = rx_engine[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:413:11  */
  assign n4504 = n4501 ? 1'b1 : n4503;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:409:9  */
  assign n4506 = n4494 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:420:27  */
  assign n4507 = rx_engine[24:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:420:35  */
  assign n4509 = n4507 == 10'b0000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:421:41  */
  assign n4510 = ctrl[15:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:422:73  */
  assign n4511 = rx_engine[14:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:422:81  */
  assign n4513 = n4511 - 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:423:50  */
  assign n4514 = rx_engine[28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:423:70  */
  assign n4515 = rx_engine[10:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:423:54  */
  assign n4516 = {n4514, n4515};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:425:73  */
  assign n4517 = rx_engine[24:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:425:82  */
  assign n4519 = n4517 - 10'b0000000001;
  assign n4520 = {n4510, n4513, n4516};
  assign n4521 = n4520[12:0]; // extract
  assign n4522 = rx_engine[14:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:420:13  */
  assign n4523 = n4509 ? n4521 : n4522;
  assign n4524 = n4520[22:13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:420:13  */
  assign n4525 = n4509 ? n4524 : n4519;
  assign n4526 = {n4525, n4523};
  assign n4527 = rx_engine[24:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:419:11  */
  assign n4528 = uart_clk ? n4526 : n4527;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:428:25  */
  assign n4529 = rx_engine[14:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:428:32  */
  assign n4531 = n4529 == 4'b0000;
  assign n4534 = rx_engine[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:428:11  */
  assign n4535 = n4531 ? 1'b0 : n4534;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:428:11  */
  assign n4536 = n4531 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:417:9  */
  assign n4538 = n4494 == 2'b11;
  assign n4540 = {n4538, n4506};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:407:7  */
  always @*
    case (n4540)
      2'b10: n4541 = n4535;
      2'b01: n4541 = n4504;
      default: n4541 = 1'b0;
    endcase
  assign n4542 = n4528[8:0]; // extract
  assign n4543 = rx_engine[10:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:407:7  */
  always @*
    case (n4540)
      2'b10: n4544 = n4542;
      2'b01: n4544 = n4543;
      default: n4544 = n4543;
    endcase
  assign n4545 = n4528[12:9]; // extract
  assign n4546 = rx_engine[14:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:407:7  */
  always @*
    case (n4540)
      2'b10: n4547 = n4545;
      2'b01: n4547 = 4'b1010;
      default: n4547 = n4546;
    endcase
  assign n4548 = n4528[22:13]; // extract
  assign n4549 = rx_engine[24:15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:407:7  */
  always @*
    case (n4540)
      2'b10: n4550 = n4548;
      2'b01: n4550 = n4497;
      default: n4550 = n4549;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:407:7  */
  always @*
    case (n4540)
      2'b10: n4551 = n4536;
      2'b01: n4551 = 1'b0;
      default: n4551 = 1'b0;
    endcase
  assign n4552 = {uart_rxd_i, n4491, n4551, n4550, n4547, n4544, n4493, n4541};
  assign n4555 = {3'b000, 1'b0, 10'b0000000000, 4'b0000, 9'b000000000, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:444:16  */
  assign n4559 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:447:16  */
  assign n4562 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:447:23  */
  assign n4563 = ~n4562;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:449:22  */
  assign n4565 = rx_fifo[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:449:45  */
  assign n4566 = rx_fifo[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:449:50  */
  assign n4567 = ~n4566;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:449:32  */
  assign n4568 = n4567 & n4565;
  assign n4570 = rx_engine[29]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:449:7  */
  assign n4571 = n4568 ? 1'b1 : n4570;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:447:7  */
  assign n4572 = n4563 ? 1'b0 : n4571;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:458:16  */
  assign n4578 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:461:16  */
  assign n4580 = ctrl[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:462:18  */
  assign n4581 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:462:25  */
  assign n4582 = ~n4581;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:463:21  */
  assign n4583 = rx_fifo[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:462:32  */
  assign n4584 = n4582 | n4583;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:462:9  */
  assign n4587 = n4584 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:461:7  */
  assign n4589 = n4580 ? n4587 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:164:5  */
  always @(posedge clk_i or posedge n4162)
    if (n4162)
      n4594 <= n4270;
    else
      n4594 <= n4264;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:324:5  */
  always @(posedge clk_i or posedge n4378)
    if (n4378)
      n4595 <= n4469;
    else
      n4595 <= n4463;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:324:5  */
  always @(posedge clk_i or posedge n4378)
    if (n4378)
      n4596 <= n4468;
    else
      n4596 <= n4462;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:316:5  */
  assign n4597 = {n4595, n4477, n4596};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:446:5  */
  always @(posedge clk_i or posedge n4559)
    if (n4559)
      n4598 <= 1'b0;
    else
      n4598 <= n4572;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:395:5  */
  always @(posedge clk_i or posedge n4481)
    if (n4481)
      n4599 <= n4555;
    else
      n4599 <= n4552;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:388:5  */
  assign n4600 = {n4598, n4599};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:444:5  */
  assign n4601 = {\rx_engine_fifo_inst.half_o , \rx_engine_fifo_inst.avail_o , \rx_engine_fifo_inst.free_o , \rx_engine_fifo_inst.rdata_o , n4345, n4354, n4346, n4343};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:316:5  */
  assign n4602 = {\tx_engine_fifo_inst.half_o , \tx_engine_fifo_inst.avail_o , \tx_engine_fifo_inst.free_o , \tx_engine_fifo_inst.rdata_o , n4295, n4308, n4302, n4293};
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:164:5  */
  always @(posedge clk_i or posedge n4162)
    if (n4162)
      n4603 <= 34'b0000000000000000000000000000000000;
    else
      n4603 <= n4265;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:460:5  */
  always @(posedge clk_i or posedge n4578)
    if (n4578)
      n4604 <= 1'b0;
    else
      n4604 <= n4589;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:303:5  */
  always @(posedge clk_i or posedge n4357)
    if (n4357)
      n4605 <= 1'b0;
    else
      n4605 <= n4372;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:262:5  */
  always @(posedge clk_i or posedge n4311)
    if (n4311)
      n4606 <= 1'b0;
    else
      n4606 <= n4323;
  /* ../../ext/neorv32/rtl/core/neorv32_uart.vhd:225:27  */
  assign n4607 = clkgen_i[n4274 * 1 +: 1]; //(Bmux)
endmodule

module neorv32_clint_1
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output [63:0] time_o,
   output mti_o,
   output msi_o);
  wire [79:0] n4062;
  wire [31:0] n4064;
  wire n4065;
  wire n4066;
  wire mtime_en;
  wire mtimecmp_en;
  wire mswi_en;
  wire [31:0] mtime_rd;
  wire [31:0] mtimecmp_rd;
  wire [31:0] mswi_rd;
  wire [63:0] mtime;
  wire ack_q;
  wire [31:0] rdata;
  wire n4070;
  wire n4071;
  wire [31:0] n4072;
  wire [31:0] neorv32_clint_mtime_inst_n4073;
  wire [63:0] neorv32_clint_mtime_inst_n4074;
  wire n4080;
  wire [12:0] n4081;
  wire n4083;
  wire n4084;
  wire n4085;
  wire n4088;
  wire [31:0] n4091;
  wire [31:0] n4096;
  wire n4097;
  wire n4098;
  wire [31:0] n4099;
  wire [31:0] neorv32_clint_mtimecmp_gen_n1_neorv32_clint_mtimecmp_inst_n4100;
  wire neorv32_clint_mtimecmp_gen_n1_neorv32_clint_mtimecmp_inst_n4101;
  wire n4107;
  wire [12:0] n4108;
  wire n4110;
  wire n4111;
  wire n4112;
  wire n4114;
  wire [31:0] n4115;
  wire [31:0] neorv32_clint_swi_gen_n1_neorv32_clint_swi_inst_n4116;
  wire neorv32_clint_swi_gen_n1_neorv32_clint_swi_inst_n4117;
  wire n4123;
  wire [13:0] n4124;
  wire n4126;
  wire n4127;
  wire n4128;
  wire [31:0] n4133;
  wire [31:0] n4135;
  wire [31:0] n4136;
  wire n4139;
  wire n4141;
  reg n4147;
  wire [33:0] n4148;
  reg [31:0] n4149;
  wire [63:0] n4150;
  assign \bus_rsp_o_bus_rsp_o[data]  = n4064; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n4065; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n4066; //(module output)
  assign time_o = n4150; //(module output)
  assign mti_o = neorv32_clint_mtimecmp_gen_n1_neorv32_clint_mtimecmp_inst_n4101; //(module output)
  assign msi_o = neorv32_clint_swi_gen_n1_neorv32_clint_swi_inst_n4117; //(module output)
  assign n4062 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n4064 = n4148[31:0]; // extract
  assign n4065 = n4148[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1026:14  */
  assign n4066 = n4148[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:86:10  */
  assign mtime_en = n4085; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:87:10  */
  assign mtimecmp_en = n4112; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:88:10  */
  assign mswi_en = n4128; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:92:10  */
  assign mtime_rd = neorv32_clint_mtime_inst_n4073; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:93:10  */
  assign mtimecmp_rd = neorv32_clint_mtimecmp_gen_n1_neorv32_clint_mtimecmp_inst_n4100; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:94:10  */
  assign mswi_rd = neorv32_clint_swi_gen_n1_neorv32_clint_swi_inst_n4116; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:97:10  */
  assign mtime = neorv32_clint_mtime_inst_n4074; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:98:10  */
  assign ack_q = n4147; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:99:10  */
  assign rdata = n4136; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:110:26  */
  assign n4070 = n4062[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:111:30  */
  assign n4071 = n4062[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:112:26  */
  assign n4072 = n4062[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:105:3  */
  neorv32_clint_mtime neorv32_clint_mtime_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .en_i(mtime_en),
    .rw_i(n4070),
    .addr_i(n4071),
    .wdata_i(n4072),
    .rdata_o(neorv32_clint_mtime_inst_n4073),
    .mtime_o(neorv32_clint_mtime_inst_n4074));
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:118:35  */
  assign n4080 = n4062[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:118:74  */
  assign n4081 = n4062[15:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:118:89  */
  assign n4083 = n4081 == 13'b1011111111111;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:118:46  */
  assign n4084 = n4083 & n4080;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:118:19  */
  assign n4085 = n4084 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:123:16  */
  assign n4088 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:126:35  */
  assign n4091 = mtime[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:130:32  */
  assign n4096 = mtime[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:143:28  */
  assign n4097 = n4062[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:144:32  */
  assign n4098 = n4062[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:145:28  */
  assign n4099 = n4062[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:138:5  */
  neorv32_clint_mtimecmp neorv32_clint_mtimecmp_gen_n1_neorv32_clint_mtimecmp_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .en_i(mtimecmp_en),
    .rw_i(n4097),
    .addr_i(n4098),
    .wdata_i(n4099),
    .mtime_i(mtime),
    .rdata_o(neorv32_clint_mtimecmp_gen_n1_neorv32_clint_mtimecmp_inst_n4100),
    .mti_o(neorv32_clint_mtimecmp_gen_n1_neorv32_clint_mtimecmp_inst_n4101));
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:152:43  */
  assign n4107 = n4062[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:152:82  */
  assign n4108 = n4062[15:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:152:97  */
  assign n4110 = n4108 == 13'b0100000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:152:54  */
  assign n4111 = n4110 & n4107;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:152:27  */
  assign n4112 = n4111 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:167:28  */
  assign n4114 = n4062[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:168:28  */
  assign n4115 = n4062[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:162:5  */
  neorv32_clint_swi neorv32_clint_swi_gen_n1_neorv32_clint_swi_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .en_i(mswi_en),
    .rw_i(n4114),
    .wdata_i(n4115),
    .rdata_o(neorv32_clint_swi_gen_n1_neorv32_clint_swi_inst_n4116),
    .swi_o(neorv32_clint_swi_gen_n1_neorv32_clint_swi_inst_n4117));
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:174:39  */
  assign n4123 = n4062[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:174:78  */
  assign n4124 = n4062[15:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:174:93  */
  assign n4126 = n4124 == 14'b00000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:174:50  */
  assign n4127 = n4126 & n4123;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:174:23  */
  assign n4128 = n4127 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:186:20  */
  assign n4133 = 32'b00000000000000000000000000000000 | mtime_rd;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:189:22  */
  assign n4135 = n4133 | mtimecmp_rd;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:193:22  */
  assign n4136 = n4135 | mswi_rd;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:204:16  */
  assign n4139 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:207:26  */
  assign n4141 = n4062[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:206:5  */
  always @(posedge clk_i or posedge n4139)
    if (n4139)
      n4147 <= 1'b0;
    else
      n4147 <= n4141;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:204:5  */
  assign n4148 = {1'b0, ack_q, rdata};
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:125:5  */
  always @(posedge clk_i or posedge n4088)
    if (n4088)
      n4149 <= 32'b00000000000000000000000000000000;
    else
      n4149 <= n4091;
  /* ../../ext/neorv32/rtl/core/neorv32_clint.vhd:123:5  */
  assign n4150 = {n4096, n4149};
endmodule

module neorv32_gpio_23
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   input  [31:0] gpio_i,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output [31:0] gpio_o,
   output cpu_irq_o);
  wire [79:0] n3228;
  wire [31:0] n3230;
  wire n3231;
  wire n3232;
  wire [22:0] port_in;
  wire [22:0] port_out;
  wire [22:0] irq_typ;
  wire [22:0] irq_pol;
  wire [22:0] irq_en;
  wire [22:0] irq_clrn;
  wire [22:0] port_in2;
  wire [22:0] irq_trig;
  wire [22:0] irq_pend;
  wire n3236;
  wire n3238;
  localparam [31:0] n3240 = 32'b00000000000000000000000000000000;
  wire n3241;
  wire n3242;
  wire [2:0] n3243;
  wire [22:0] n3244;
  wire n3246;
  wire [22:0] n3247;
  wire n3249;
  wire [22:0] n3250;
  wire n3252;
  wire [22:0] n3253;
  wire n3255;
  wire [22:0] n3256;
  wire n3258;
  wire [4:0] n3259;
  reg [22:0] n3260;
  reg [22:0] n3261;
  reg [22:0] n3262;
  reg [22:0] n3263;
  reg [22:0] n3265;
  wire [2:0] n3266;
  wire n3268;
  wire n3270;
  wire n3272;
  wire n3274;
  wire n3276;
  wire n3278;
  wire [5:0] n3279;
  wire [22:0] n3280;
  reg [22:0] n3281;
  wire [22:0] n3282;
  wire [22:0] n3283;
  wire [22:0] n3289;
  wire [22:0] n3290;
  wire [22:0] n3291;
  wire [8:0] n3292;
  wire n3293;
  wire n3294;
  wire n3295;
  wire n3296;
  wire [22:0] n3298;
  wire [33:0] n3300;
  wire n3321;
  wire [22:0] n3323;
  localparam [31:0] n3332 = 32'b00000000000000000000000000000000;
  wire [8:0] n3333;
  wire n3337;
  wire n3338;
  wire [1:0] n3339;
  wire n3340;
  wire n3341;
  wire n3343;
  wire n3344;
  wire n3346;
  wire n3347;
  wire n3348;
  wire n3349;
  wire n3350;
  wire n3352;
  wire n3353;
  wire n3354;
  wire n3355;
  wire n3356;
  wire n3358;
  wire [3:0] n3360;
  reg n3361;
  wire n3365;
  wire n3366;
  wire [1:0] n3367;
  wire n3368;
  wire n3369;
  wire n3371;
  wire n3372;
  wire n3374;
  wire n3375;
  wire n3376;
  wire n3377;
  wire n3378;
  wire n3380;
  wire n3381;
  wire n3382;
  wire n3383;
  wire n3384;
  wire n3386;
  wire [3:0] n3388;
  reg n3389;
  wire n3393;
  wire n3394;
  wire [1:0] n3395;
  wire n3396;
  wire n3397;
  wire n3399;
  wire n3400;
  wire n3402;
  wire n3403;
  wire n3404;
  wire n3405;
  wire n3406;
  wire n3408;
  wire n3409;
  wire n3410;
  wire n3411;
  wire n3412;
  wire n3414;
  wire [3:0] n3416;
  reg n3417;
  wire n3421;
  wire n3422;
  wire [1:0] n3423;
  wire n3424;
  wire n3425;
  wire n3427;
  wire n3428;
  wire n3430;
  wire n3431;
  wire n3432;
  wire n3433;
  wire n3434;
  wire n3436;
  wire n3437;
  wire n3438;
  wire n3439;
  wire n3440;
  wire n3442;
  wire [3:0] n3444;
  reg n3445;
  wire n3449;
  wire n3450;
  wire [1:0] n3451;
  wire n3452;
  wire n3453;
  wire n3455;
  wire n3456;
  wire n3458;
  wire n3459;
  wire n3460;
  wire n3461;
  wire n3462;
  wire n3464;
  wire n3465;
  wire n3466;
  wire n3467;
  wire n3468;
  wire n3470;
  wire [3:0] n3472;
  reg n3473;
  wire n3477;
  wire n3478;
  wire [1:0] n3479;
  wire n3480;
  wire n3481;
  wire n3483;
  wire n3484;
  wire n3486;
  wire n3487;
  wire n3488;
  wire n3489;
  wire n3490;
  wire n3492;
  wire n3493;
  wire n3494;
  wire n3495;
  wire n3496;
  wire n3498;
  wire [3:0] n3500;
  reg n3501;
  wire n3505;
  wire n3506;
  wire [1:0] n3507;
  wire n3508;
  wire n3509;
  wire n3511;
  wire n3512;
  wire n3514;
  wire n3515;
  wire n3516;
  wire n3517;
  wire n3518;
  wire n3520;
  wire n3521;
  wire n3522;
  wire n3523;
  wire n3524;
  wire n3526;
  wire [3:0] n3528;
  reg n3529;
  wire n3533;
  wire n3534;
  wire [1:0] n3535;
  wire n3536;
  wire n3537;
  wire n3539;
  wire n3540;
  wire n3542;
  wire n3543;
  wire n3544;
  wire n3545;
  wire n3546;
  wire n3548;
  wire n3549;
  wire n3550;
  wire n3551;
  wire n3552;
  wire n3554;
  wire [3:0] n3556;
  reg n3557;
  wire n3561;
  wire n3562;
  wire [1:0] n3563;
  wire n3564;
  wire n3565;
  wire n3567;
  wire n3568;
  wire n3570;
  wire n3571;
  wire n3572;
  wire n3573;
  wire n3574;
  wire n3576;
  wire n3577;
  wire n3578;
  wire n3579;
  wire n3580;
  wire n3582;
  wire [3:0] n3584;
  reg n3585;
  wire n3589;
  wire n3590;
  wire [1:0] n3591;
  wire n3592;
  wire n3593;
  wire n3595;
  wire n3596;
  wire n3598;
  wire n3599;
  wire n3600;
  wire n3601;
  wire n3602;
  wire n3604;
  wire n3605;
  wire n3606;
  wire n3607;
  wire n3608;
  wire n3610;
  wire [3:0] n3612;
  reg n3613;
  wire n3617;
  wire n3618;
  wire [1:0] n3619;
  wire n3620;
  wire n3621;
  wire n3623;
  wire n3624;
  wire n3626;
  wire n3627;
  wire n3628;
  wire n3629;
  wire n3630;
  wire n3632;
  wire n3633;
  wire n3634;
  wire n3635;
  wire n3636;
  wire n3638;
  wire [3:0] n3640;
  reg n3641;
  wire n3645;
  wire n3646;
  wire [1:0] n3647;
  wire n3648;
  wire n3649;
  wire n3651;
  wire n3652;
  wire n3654;
  wire n3655;
  wire n3656;
  wire n3657;
  wire n3658;
  wire n3660;
  wire n3661;
  wire n3662;
  wire n3663;
  wire n3664;
  wire n3666;
  wire [3:0] n3668;
  reg n3669;
  wire n3673;
  wire n3674;
  wire [1:0] n3675;
  wire n3676;
  wire n3677;
  wire n3679;
  wire n3680;
  wire n3682;
  wire n3683;
  wire n3684;
  wire n3685;
  wire n3686;
  wire n3688;
  wire n3689;
  wire n3690;
  wire n3691;
  wire n3692;
  wire n3694;
  wire [3:0] n3696;
  reg n3697;
  wire n3701;
  wire n3702;
  wire [1:0] n3703;
  wire n3704;
  wire n3705;
  wire n3707;
  wire n3708;
  wire n3710;
  wire n3711;
  wire n3712;
  wire n3713;
  wire n3714;
  wire n3716;
  wire n3717;
  wire n3718;
  wire n3719;
  wire n3720;
  wire n3722;
  wire [3:0] n3724;
  reg n3725;
  wire n3729;
  wire n3730;
  wire [1:0] n3731;
  wire n3732;
  wire n3733;
  wire n3735;
  wire n3736;
  wire n3738;
  wire n3739;
  wire n3740;
  wire n3741;
  wire n3742;
  wire n3744;
  wire n3745;
  wire n3746;
  wire n3747;
  wire n3748;
  wire n3750;
  wire [3:0] n3752;
  reg n3753;
  wire n3757;
  wire n3758;
  wire [1:0] n3759;
  wire n3760;
  wire n3761;
  wire n3763;
  wire n3764;
  wire n3766;
  wire n3767;
  wire n3768;
  wire n3769;
  wire n3770;
  wire n3772;
  wire n3773;
  wire n3774;
  wire n3775;
  wire n3776;
  wire n3778;
  wire [3:0] n3780;
  reg n3781;
  wire n3785;
  wire n3786;
  wire [1:0] n3787;
  wire n3788;
  wire n3789;
  wire n3791;
  wire n3792;
  wire n3794;
  wire n3795;
  wire n3796;
  wire n3797;
  wire n3798;
  wire n3800;
  wire n3801;
  wire n3802;
  wire n3803;
  wire n3804;
  wire n3806;
  wire [3:0] n3808;
  reg n3809;
  wire n3813;
  wire n3814;
  wire [1:0] n3815;
  wire n3816;
  wire n3817;
  wire n3819;
  wire n3820;
  wire n3822;
  wire n3823;
  wire n3824;
  wire n3825;
  wire n3826;
  wire n3828;
  wire n3829;
  wire n3830;
  wire n3831;
  wire n3832;
  wire n3834;
  wire [3:0] n3836;
  reg n3837;
  wire n3841;
  wire n3842;
  wire [1:0] n3843;
  wire n3844;
  wire n3845;
  wire n3847;
  wire n3848;
  wire n3850;
  wire n3851;
  wire n3852;
  wire n3853;
  wire n3854;
  wire n3856;
  wire n3857;
  wire n3858;
  wire n3859;
  wire n3860;
  wire n3862;
  wire [3:0] n3864;
  reg n3865;
  wire n3869;
  wire n3870;
  wire [1:0] n3871;
  wire n3872;
  wire n3873;
  wire n3875;
  wire n3876;
  wire n3878;
  wire n3879;
  wire n3880;
  wire n3881;
  wire n3882;
  wire n3884;
  wire n3885;
  wire n3886;
  wire n3887;
  wire n3888;
  wire n3890;
  wire [3:0] n3892;
  reg n3893;
  wire n3897;
  wire n3898;
  wire [1:0] n3899;
  wire n3900;
  wire n3901;
  wire n3903;
  wire n3904;
  wire n3906;
  wire n3907;
  wire n3908;
  wire n3909;
  wire n3910;
  wire n3912;
  wire n3913;
  wire n3914;
  wire n3915;
  wire n3916;
  wire n3918;
  wire [3:0] n3920;
  reg n3921;
  wire n3925;
  wire n3926;
  wire [1:0] n3927;
  wire n3928;
  wire n3929;
  wire n3931;
  wire n3932;
  wire n3934;
  wire n3935;
  wire n3936;
  wire n3937;
  wire n3938;
  wire n3940;
  wire n3941;
  wire n3942;
  wire n3943;
  wire n3944;
  wire n3946;
  wire [3:0] n3948;
  reg n3949;
  wire n3953;
  wire n3954;
  wire [1:0] n3955;
  wire n3956;
  wire n3957;
  wire n3959;
  wire n3960;
  wire n3962;
  wire n3963;
  wire n3964;
  wire n3965;
  wire n3966;
  wire n3968;
  wire n3969;
  wire n3970;
  wire n3971;
  wire n3972;
  wire n3974;
  wire [3:0] n3976;
  reg n3977;
  wire n3980;
  wire [22:0] n3982;
  wire [22:0] n3983;
  wire [22:0] n3984;
  wire n3991;
  wire n3993;
  wire n3995;
  wire n3996;
  wire n3997;
  wire n3998;
  wire n3999;
  wire n4000;
  wire n4001;
  wire n4002;
  wire n4003;
  wire n4004;
  wire n4005;
  wire n4006;
  wire n4007;
  wire n4008;
  wire n4009;
  wire n4010;
  wire n4011;
  wire n4012;
  wire n4013;
  wire n4014;
  wire n4015;
  wire n4016;
  wire n4017;
  wire n4018;
  wire n4019;
  wire n4020;
  wire n4021;
  wire n4022;
  wire n4023;
  wire n4024;
  wire n4025;
  wire n4026;
  wire n4027;
  wire n4028;
  wire n4029;
  wire n4030;
  wire n4031;
  wire n4032;
  wire n4033;
  wire n4034;
  wire n4035;
  wire n4036;
  wire n4037;
  wire n4038;
  reg [22:0] n4046;
  wire [22:0] n4047;
  reg [22:0] n4048;
  wire [22:0] n4049;
  reg [22:0] n4050;
  wire [22:0] n4051;
  reg [22:0] n4052;
  wire [22:0] n4053;
  reg [22:0] n4054;
  reg [22:0] n4055;
  reg [22:0] n4056;
  wire [22:0] n4057;
  reg [22:0] n4058;
  reg [33:0] n4059;
  wire [31:0] n4060;
  reg n4061;
  assign \bus_rsp_o_bus_rsp_o[data]  = n3230; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n3231; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n3232; //(module output)
  assign gpio_o = n4060; //(module output)
  assign cpu_irq_o = n4061; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:48:25  */
  assign n3228 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n3230 = n4059[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:55:3  */
  assign n3231 = n4059[32]; // extract
  assign n3232 = n4059[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:44:10  */
  assign port_in = n4046; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:44:19  */
  assign port_out = n4048; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:45:10  */
  assign irq_typ = n4050; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:45:19  */
  assign irq_pol = n4052; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:46:10  */
  assign irq_en = n4054; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:46:18  */
  assign irq_clrn = n4055; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:49:10  */
  assign port_in2 = n4056; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:49:20  */
  assign irq_trig = n4057; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:49:30  */
  assign irq_pend = n4058; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:57:16  */
  assign n3236 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:66:35  */
  assign n3238 = n3228[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:71:21  */
  assign n3241 = n3228[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:72:23  */
  assign n3242 = n3228[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:73:30  */
  assign n3243 = n3228[4:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:74:58  */
  assign n3244 = n3228[54:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:74:13  */
  assign n3246 = n3243 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:75:58  */
  assign n3247 = n3228[54:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:75:13  */
  assign n3249 = n3243 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:76:58  */
  assign n3250 = n3228[54:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:76:13  */
  assign n3252 = n3243 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:77:58  */
  assign n3253 = n3228[54:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:77:13  */
  assign n3255 = n3243 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:78:58  */
  assign n3256 = n3228[54:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:78:13  */
  assign n3258 = n3243 == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:44  */
  assign n3259 = {n3258, n3255, n3252, n3249, n3246};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:73:11  */
  always @*
    case (n3259)
      5'b10000: n3260 = port_out;
      5'b01000: n3260 = port_out;
      5'b00100: n3260 = port_out;
      5'b00010: n3260 = port_out;
      5'b00001: n3260 = n3244;
      default: n3260 = port_out;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:73:11  */
  always @*
    case (n3259)
      5'b10000: n3261 = irq_typ;
      5'b01000: n3261 = irq_typ;
      5'b00100: n3261 = irq_typ;
      5'b00010: n3261 = n3247;
      5'b00001: n3261 = irq_typ;
      default: n3261 = irq_typ;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:73:11  */
  always @*
    case (n3259)
      5'b10000: n3262 = irq_pol;
      5'b01000: n3262 = irq_pol;
      5'b00100: n3262 = n3250;
      5'b00010: n3262 = irq_pol;
      5'b00001: n3262 = irq_pol;
      default: n3262 = irq_pol;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:73:11  */
  always @*
    case (n3259)
      5'b10000: n3263 = irq_en;
      5'b01000: n3263 = n3253;
      5'b00100: n3263 = irq_en;
      5'b00010: n3263 = irq_en;
      5'b00001: n3263 = irq_en;
      default: n3263 = irq_en;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:73:11  */
  always @*
    case (n3259)
      5'b10000: n3265 = n3256;
      5'b01000: n3265 = 23'b11111111111111111111111;
      5'b00100: n3265 = 23'b11111111111111111111111;
      5'b00010: n3265 = 23'b11111111111111111111111;
      5'b00001: n3265 = 23'b11111111111111111111111;
      default: n3265 = 23'b11111111111111111111111;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:82:30  */
  assign n3266 = n3228[4:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:83:13  */
  assign n3268 = n3266 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:84:13  */
  assign n3270 = n3266 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:85:13  */
  assign n3272 = n3266 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:86:13  */
  assign n3274 = n3266 == 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:87:13  */
  assign n3276 = n3266 == 3'b110;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:88:13  */
  assign n3278 = n3266 == 3'b111;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:702:7  */
  assign n3279 = {n3278, n3276, n3274, n3272, n3270, n3268};
  assign n3280 = n3240[22:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:82:11  */
  always @*
    case (n3279)
      6'b100000: n3281 = irq_pend;
      6'b010000: n3281 = irq_en;
      6'b001000: n3281 = irq_pol;
      6'b000100: n3281 = irq_typ;
      6'b000010: n3281 = port_out;
      6'b000001: n3281 = port_in;
      default: n3281 = n3280;
    endcase
  assign n3282 = n3240[22:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:72:9  */
  assign n3283 = n3242 ? n3282 : n3281;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:72:9  */
  assign n3289 = n3242 ? n3265 : 23'b11111111111111111111111;
  assign n3290 = n3240[22:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:71:7  */
  assign n3291 = n3241 ? n3283 : n3290;
  assign n3292 = n3240[31:23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:71:7  */
  assign n3293 = n3242 & n3241;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:71:7  */
  assign n3294 = n3242 & n3241;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:71:7  */
  assign n3295 = n3242 & n3241;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:71:7  */
  assign n3296 = n3242 & n3241;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:71:7  */
  assign n3298 = n3241 ? n3289 : 23'b11111111111111111111111;
  assign n3300 = {1'b0, n3238, n3292, n3291};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:99:16  */
  assign n3321 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:103:25  */
  assign n3323 = gpio_i[22:0]; // extract
  assign n3333 = n3332[31:23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3337 = irq_typ[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3338 = irq_pol[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3339 = {n3337, n3338};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3340 = port_in[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3341 = ~n3340;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3343 = n3339 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3344 = port_in[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3346 = n3339 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3347 = port_in[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3348 = ~n3347;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3349 = port_in2[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3350 = n3348 & n3349;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3352 = n3339 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3353 = port_in[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3354 = port_in2[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3355 = ~n3354;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3356 = n3353 & n3355;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3358 = n3339 == 2'b11;
  assign n3360 = {n3358, n3352, n3346, n3343};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3360)
      4'b1000: n3361 = n3356;
      4'b0100: n3361 = n3350;
      4'b0010: n3361 = n3344;
      4'b0001: n3361 = n3341;
      default: n3361 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3365 = irq_typ[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3366 = irq_pol[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3367 = {n3365, n3366};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3368 = port_in[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3369 = ~n3368;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3371 = n3367 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3372 = port_in[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3374 = n3367 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3375 = port_in[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3376 = ~n3375;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3377 = port_in2[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3378 = n3376 & n3377;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3380 = n3367 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3381 = port_in[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3382 = port_in2[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3383 = ~n3382;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3384 = n3381 & n3383;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3386 = n3367 == 2'b11;
  assign n3388 = {n3386, n3380, n3374, n3371};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3388)
      4'b1000: n3389 = n3384;
      4'b0100: n3389 = n3378;
      4'b0010: n3389 = n3372;
      4'b0001: n3389 = n3369;
      default: n3389 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3393 = irq_typ[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3394 = irq_pol[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3395 = {n3393, n3394};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3396 = port_in[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3397 = ~n3396;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3399 = n3395 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3400 = port_in[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3402 = n3395 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3403 = port_in[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3404 = ~n3403;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3405 = port_in2[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3406 = n3404 & n3405;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3408 = n3395 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3409 = port_in[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3410 = port_in2[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3411 = ~n3410;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3412 = n3409 & n3411;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3414 = n3395 == 2'b11;
  assign n3416 = {n3414, n3408, n3402, n3399};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3416)
      4'b1000: n3417 = n3412;
      4'b0100: n3417 = n3406;
      4'b0010: n3417 = n3400;
      4'b0001: n3417 = n3397;
      default: n3417 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3421 = irq_typ[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3422 = irq_pol[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3423 = {n3421, n3422};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3424 = port_in[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3425 = ~n3424;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3427 = n3423 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3428 = port_in[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3430 = n3423 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3431 = port_in[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3432 = ~n3431;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3433 = port_in2[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3434 = n3432 & n3433;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3436 = n3423 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3437 = port_in[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3438 = port_in2[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3439 = ~n3438;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3440 = n3437 & n3439;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3442 = n3423 == 2'b11;
  assign n3444 = {n3442, n3436, n3430, n3427};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3444)
      4'b1000: n3445 = n3440;
      4'b0100: n3445 = n3434;
      4'b0010: n3445 = n3428;
      4'b0001: n3445 = n3425;
      default: n3445 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3449 = irq_typ[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3450 = irq_pol[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3451 = {n3449, n3450};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3452 = port_in[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3453 = ~n3452;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3455 = n3451 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3456 = port_in[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3458 = n3451 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3459 = port_in[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3460 = ~n3459;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3461 = port_in2[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3462 = n3460 & n3461;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3464 = n3451 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3465 = port_in[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3466 = port_in2[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3467 = ~n3466;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3468 = n3465 & n3467;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3470 = n3451 == 2'b11;
  assign n3472 = {n3470, n3464, n3458, n3455};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3472)
      4'b1000: n3473 = n3468;
      4'b0100: n3473 = n3462;
      4'b0010: n3473 = n3456;
      4'b0001: n3473 = n3453;
      default: n3473 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3477 = irq_typ[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3478 = irq_pol[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3479 = {n3477, n3478};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3480 = port_in[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3481 = ~n3480;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3483 = n3479 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3484 = port_in[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3486 = n3479 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3487 = port_in[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3488 = ~n3487;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3489 = port_in2[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3490 = n3488 & n3489;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3492 = n3479 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3493 = port_in[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3494 = port_in2[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3495 = ~n3494;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3496 = n3493 & n3495;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3498 = n3479 == 2'b11;
  assign n3500 = {n3498, n3492, n3486, n3483};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3500)
      4'b1000: n3501 = n3496;
      4'b0100: n3501 = n3490;
      4'b0010: n3501 = n3484;
      4'b0001: n3501 = n3481;
      default: n3501 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3505 = irq_typ[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3506 = irq_pol[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3507 = {n3505, n3506};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3508 = port_in[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3509 = ~n3508;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3511 = n3507 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3512 = port_in[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3514 = n3507 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3515 = port_in[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3516 = ~n3515;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3517 = port_in2[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3518 = n3516 & n3517;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3520 = n3507 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3521 = port_in[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3522 = port_in2[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3523 = ~n3522;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3524 = n3521 & n3523;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3526 = n3507 == 2'b11;
  assign n3528 = {n3526, n3520, n3514, n3511};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3528)
      4'b1000: n3529 = n3524;
      4'b0100: n3529 = n3518;
      4'b0010: n3529 = n3512;
      4'b0001: n3529 = n3509;
      default: n3529 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3533 = irq_typ[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3534 = irq_pol[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3535 = {n3533, n3534};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3536 = port_in[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3537 = ~n3536;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3539 = n3535 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3540 = port_in[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3542 = n3535 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3543 = port_in[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3544 = ~n3543;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3545 = port_in2[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3546 = n3544 & n3545;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3548 = n3535 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3549 = port_in[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3550 = port_in2[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3551 = ~n3550;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3552 = n3549 & n3551;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3554 = n3535 == 2'b11;
  assign n3556 = {n3554, n3548, n3542, n3539};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3556)
      4'b1000: n3557 = n3552;
      4'b0100: n3557 = n3546;
      4'b0010: n3557 = n3540;
      4'b0001: n3557 = n3537;
      default: n3557 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3561 = irq_typ[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3562 = irq_pol[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3563 = {n3561, n3562};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3564 = port_in[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3565 = ~n3564;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3567 = n3563 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3568 = port_in[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3570 = n3563 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3571 = port_in[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3572 = ~n3571;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3573 = port_in2[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3574 = n3572 & n3573;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3576 = n3563 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3577 = port_in[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3578 = port_in2[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3579 = ~n3578;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3580 = n3577 & n3579;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3582 = n3563 == 2'b11;
  assign n3584 = {n3582, n3576, n3570, n3567};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3584)
      4'b1000: n3585 = n3580;
      4'b0100: n3585 = n3574;
      4'b0010: n3585 = n3568;
      4'b0001: n3585 = n3565;
      default: n3585 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3589 = irq_typ[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3590 = irq_pol[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3591 = {n3589, n3590};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3592 = port_in[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3593 = ~n3592;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3595 = n3591 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3596 = port_in[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3598 = n3591 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3599 = port_in[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3600 = ~n3599;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3601 = port_in2[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3602 = n3600 & n3601;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3604 = n3591 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3605 = port_in[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3606 = port_in2[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3607 = ~n3606;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3608 = n3605 & n3607;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3610 = n3591 == 2'b11;
  assign n3612 = {n3610, n3604, n3598, n3595};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3612)
      4'b1000: n3613 = n3608;
      4'b0100: n3613 = n3602;
      4'b0010: n3613 = n3596;
      4'b0001: n3613 = n3593;
      default: n3613 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3617 = irq_typ[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3618 = irq_pol[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3619 = {n3617, n3618};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3620 = port_in[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3621 = ~n3620;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3623 = n3619 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3624 = port_in[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3626 = n3619 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3627 = port_in[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3628 = ~n3627;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3629 = port_in2[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3630 = n3628 & n3629;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3632 = n3619 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3633 = port_in[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3634 = port_in2[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3635 = ~n3634;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3636 = n3633 & n3635;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3638 = n3619 == 2'b11;
  assign n3640 = {n3638, n3632, n3626, n3623};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3640)
      4'b1000: n3641 = n3636;
      4'b0100: n3641 = n3630;
      4'b0010: n3641 = n3624;
      4'b0001: n3641 = n3621;
      default: n3641 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3645 = irq_typ[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3646 = irq_pol[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3647 = {n3645, n3646};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3648 = port_in[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3649 = ~n3648;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3651 = n3647 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3652 = port_in[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3654 = n3647 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3655 = port_in[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3656 = ~n3655;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3657 = port_in2[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3658 = n3656 & n3657;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3660 = n3647 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3661 = port_in[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3662 = port_in2[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3663 = ~n3662;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3664 = n3661 & n3663;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3666 = n3647 == 2'b11;
  assign n3668 = {n3666, n3660, n3654, n3651};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3668)
      4'b1000: n3669 = n3664;
      4'b0100: n3669 = n3658;
      4'b0010: n3669 = n3652;
      4'b0001: n3669 = n3649;
      default: n3669 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3673 = irq_typ[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3674 = irq_pol[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3675 = {n3673, n3674};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3676 = port_in[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3677 = ~n3676;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3679 = n3675 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3680 = port_in[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3682 = n3675 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3683 = port_in[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3684 = ~n3683;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3685 = port_in2[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3686 = n3684 & n3685;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3688 = n3675 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3689 = port_in[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3690 = port_in2[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3691 = ~n3690;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3692 = n3689 & n3691;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3694 = n3675 == 2'b11;
  assign n3696 = {n3694, n3688, n3682, n3679};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3696)
      4'b1000: n3697 = n3692;
      4'b0100: n3697 = n3686;
      4'b0010: n3697 = n3680;
      4'b0001: n3697 = n3677;
      default: n3697 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3701 = irq_typ[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3702 = irq_pol[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3703 = {n3701, n3702};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3704 = port_in[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3705 = ~n3704;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3707 = n3703 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3708 = port_in[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3710 = n3703 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3711 = port_in[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3712 = ~n3711;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3713 = port_in2[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3714 = n3712 & n3713;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3716 = n3703 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3717 = port_in[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3718 = port_in2[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3719 = ~n3718;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3720 = n3717 & n3719;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3722 = n3703 == 2'b11;
  assign n3724 = {n3722, n3716, n3710, n3707};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3724)
      4'b1000: n3725 = n3720;
      4'b0100: n3725 = n3714;
      4'b0010: n3725 = n3708;
      4'b0001: n3725 = n3705;
      default: n3725 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3729 = irq_typ[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3730 = irq_pol[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3731 = {n3729, n3730};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3732 = port_in[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3733 = ~n3732;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3735 = n3731 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3736 = port_in[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3738 = n3731 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3739 = port_in[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3740 = ~n3739;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3741 = port_in2[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3742 = n3740 & n3741;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3744 = n3731 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3745 = port_in[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3746 = port_in2[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3747 = ~n3746;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3748 = n3745 & n3747;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3750 = n3731 == 2'b11;
  assign n3752 = {n3750, n3744, n3738, n3735};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3752)
      4'b1000: n3753 = n3748;
      4'b0100: n3753 = n3742;
      4'b0010: n3753 = n3736;
      4'b0001: n3753 = n3733;
      default: n3753 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3757 = irq_typ[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3758 = irq_pol[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3759 = {n3757, n3758};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3760 = port_in[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3761 = ~n3760;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3763 = n3759 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3764 = port_in[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3766 = n3759 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3767 = port_in[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3768 = ~n3767;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3769 = port_in2[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3770 = n3768 & n3769;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3772 = n3759 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3773 = port_in[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3774 = port_in2[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3775 = ~n3774;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3776 = n3773 & n3775;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3778 = n3759 == 2'b11;
  assign n3780 = {n3778, n3772, n3766, n3763};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3780)
      4'b1000: n3781 = n3776;
      4'b0100: n3781 = n3770;
      4'b0010: n3781 = n3764;
      4'b0001: n3781 = n3761;
      default: n3781 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3785 = irq_typ[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3786 = irq_pol[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3787 = {n3785, n3786};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3788 = port_in[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3789 = ~n3788;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3791 = n3787 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3792 = port_in[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3794 = n3787 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3795 = port_in[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3796 = ~n3795;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3797 = port_in2[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3798 = n3796 & n3797;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3800 = n3787 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3801 = port_in[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3802 = port_in2[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3803 = ~n3802;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3804 = n3801 & n3803;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3806 = n3787 == 2'b11;
  assign n3808 = {n3806, n3800, n3794, n3791};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3808)
      4'b1000: n3809 = n3804;
      4'b0100: n3809 = n3798;
      4'b0010: n3809 = n3792;
      4'b0001: n3809 = n3789;
      default: n3809 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3813 = irq_typ[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3814 = irq_pol[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3815 = {n3813, n3814};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3816 = port_in[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3817 = ~n3816;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3819 = n3815 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3820 = port_in[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3822 = n3815 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3823 = port_in[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3824 = ~n3823;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3825 = port_in2[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3826 = n3824 & n3825;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3828 = n3815 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3829 = port_in[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3830 = port_in2[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3831 = ~n3830;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3832 = n3829 & n3831;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3834 = n3815 == 2'b11;
  assign n3836 = {n3834, n3828, n3822, n3819};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3836)
      4'b1000: n3837 = n3832;
      4'b0100: n3837 = n3826;
      4'b0010: n3837 = n3820;
      4'b0001: n3837 = n3817;
      default: n3837 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3841 = irq_typ[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3842 = irq_pol[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3843 = {n3841, n3842};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3844 = port_in[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3845 = ~n3844;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3847 = n3843 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3848 = port_in[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3850 = n3843 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3851 = port_in[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3852 = ~n3851;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3853 = port_in2[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3854 = n3852 & n3853;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3856 = n3843 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3857 = port_in[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3858 = port_in2[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3859 = ~n3858;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3860 = n3857 & n3859;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3862 = n3843 == 2'b11;
  assign n3864 = {n3862, n3856, n3850, n3847};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3864)
      4'b1000: n3865 = n3860;
      4'b0100: n3865 = n3854;
      4'b0010: n3865 = n3848;
      4'b0001: n3865 = n3845;
      default: n3865 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3869 = irq_typ[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3870 = irq_pol[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3871 = {n3869, n3870};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3872 = port_in[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3873 = ~n3872;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3875 = n3871 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3876 = port_in[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3878 = n3871 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3879 = port_in[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3880 = ~n3879;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3881 = port_in2[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3882 = n3880 & n3881;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3884 = n3871 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3885 = port_in[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3886 = port_in2[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3887 = ~n3886;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3888 = n3885 & n3887;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3890 = n3871 == 2'b11;
  assign n3892 = {n3890, n3884, n3878, n3875};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3892)
      4'b1000: n3893 = n3888;
      4'b0100: n3893 = n3882;
      4'b0010: n3893 = n3876;
      4'b0001: n3893 = n3873;
      default: n3893 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3897 = irq_typ[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3898 = irq_pol[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3899 = {n3897, n3898};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3900 = port_in[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3901 = ~n3900;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3903 = n3899 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3904 = port_in[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3906 = n3899 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3907 = port_in[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3908 = ~n3907;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3909 = port_in2[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3910 = n3908 & n3909;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3912 = n3899 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3913 = port_in[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3914 = port_in2[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3915 = ~n3914;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3916 = n3913 & n3915;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3918 = n3899 == 2'b11;
  assign n3920 = {n3918, n3912, n3906, n3903};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3920)
      4'b1000: n3921 = n3916;
      4'b0100: n3921 = n3910;
      4'b0010: n3921 = n3904;
      4'b0001: n3921 = n3901;
      default: n3921 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3925 = irq_typ[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3926 = irq_pol[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3927 = {n3925, n3926};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3928 = port_in[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3929 = ~n3928;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3931 = n3927 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3932 = port_in[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3934 = n3927 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3935 = port_in[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3936 = ~n3935;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3937 = port_in2[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3938 = n3936 & n3937;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3940 = n3927 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3941 = port_in[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3942 = port_in2[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3943 = ~n3942;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3944 = n3941 & n3943;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3946 = n3927 == 2'b11;
  assign n3948 = {n3946, n3940, n3934, n3931};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3948)
      4'b1000: n3949 = n3944;
      4'b0100: n3949 = n3938;
      4'b0010: n3949 = n3932;
      4'b0001: n3949 = n3929;
      default: n3949 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:23  */
  assign n3953 = irq_typ[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:36  */
  assign n3954 = irq_pol[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:123:27  */
  assign n3955 = {n3953, n3954};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:50  */
  assign n3956 = port_in[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:39  */
  assign n3957 = ~n3956;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:125:9  */
  assign n3959 = n3955 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:46  */
  assign n3960 = port_in[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:126:9  */
  assign n3962 = n3955 == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:51  */
  assign n3963 = port_in[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:40  */
  assign n3964 = ~n3963;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:68  */
  assign n3965 = port_in2[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:56  */
  assign n3966 = n3964 & n3965;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:127:9  */
  assign n3968 = n3955 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:46  */
  assign n3969 = port_in[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:67  */
  assign n3970 = port_in2[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:55  */
  assign n3971 = ~n3970;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:50  */
  assign n3972 = n3969 & n3971;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:128:9  */
  assign n3974 = n3955 == 2'b11;
  assign n3976 = {n3974, n3968, n3962, n3959};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:124:7  */
  always @*
    case (n3976)
      4'b1000: n3977 = n3972;
      4'b0100: n3977 = n3966;
      4'b0010: n3977 = n3960;
      4'b0001: n3977 = n3957;
      default: n3977 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:137:16  */
  assign n3980 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:141:42  */
  assign n3982 = irq_pend & irq_clrn;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:141:56  */
  assign n3983 = n3982 | irq_trig;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:141:27  */
  assign n3984 = irq_en & n3983;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n3991 = irq_pend[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n3993 = 1'b0 | n3991;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n3995 = irq_pend[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n3996 = n3993 | n3995;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n3997 = irq_pend[20]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n3998 = n3996 | n3997;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n3999 = irq_pend[19]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4000 = n3998 | n3999;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4001 = irq_pend[18]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4002 = n4000 | n4001;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4003 = irq_pend[17]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4004 = n4002 | n4003;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4005 = irq_pend[16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4006 = n4004 | n4005;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4007 = irq_pend[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4008 = n4006 | n4007;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4009 = irq_pend[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4010 = n4008 | n4009;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4011 = irq_pend[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4012 = n4010 | n4011;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4013 = irq_pend[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4014 = n4012 | n4013;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4015 = irq_pend[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4016 = n4014 | n4015;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4017 = irq_pend[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4018 = n4016 | n4017;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4019 = irq_pend[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4020 = n4018 | n4019;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4021 = irq_pend[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4022 = n4020 | n4021;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4023 = irq_pend[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4024 = n4022 | n4023;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4025 = irq_pend[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4026 = n4024 | n4025;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4027 = irq_pend[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4028 = n4026 | n4027;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4029 = irq_pend[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4030 = n4028 | n4029;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4031 = irq_pend[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4032 = n4030 | n4031;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4033 = irq_pend[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4034 = n4032 | n4033;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4035 = irq_pend[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4036 = n4034 | n4035;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n4037 = irq_pend[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n4038 = n4036 | n4037;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:102:5  */
  always @(posedge clk_i or posedge n3321)
    if (n3321)
      n4046 <= 23'b00000000000000000000000;
    else
      n4046 <= n3323;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  assign n4047 = n3293 ? n3260 : port_out;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  always @(posedge clk_i or posedge n3236)
    if (n3236)
      n4048 <= 23'b00000000000000000000000;
    else
      n4048 <= n4047;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  assign n4049 = n3294 ? n3261 : irq_typ;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  always @(posedge clk_i or posedge n3236)
    if (n3236)
      n4050 <= 23'b00000000000000000000000;
    else
      n4050 <= n4049;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  assign n4051 = n3295 ? n3262 : irq_pol;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  always @(posedge clk_i or posedge n3236)
    if (n3236)
      n4052 <= 23'b00000000000000000000000;
    else
      n4052 <= n4051;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  assign n4053 = n3296 ? n3263 : irq_en;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  always @(posedge clk_i or posedge n3236)
    if (n3236)
      n4054 <= 23'b00000000000000000000000;
    else
      n4054 <= n4053;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  always @(posedge clk_i or posedge n3236)
    if (n3236)
      n4055 <= 23'b00000000000000000000000;
    else
      n4055 <= n3298;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:102:5  */
  always @(posedge clk_i or posedge n3321)
    if (n3321)
      n4056 <= 23'b00000000000000000000000;
    else
      n4056 <= port_in;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:99:5  */
  assign n4057 = {n3977, n3949, n3921, n3893, n3865, n3837, n3809, n3781, n3753, n3725, n3697, n3669, n3641, n3613, n3585, n3557, n3529, n3501, n3473, n3445, n3417, n3389, n3361};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:140:5  */
  always @(posedge clk_i or posedge n3980)
    if (n3980)
      n4058 <= 23'b00000000000000000000000;
    else
      n4058 <= n3984;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:64:5  */
  always @(posedge clk_i or posedge n3236)
    if (n3236)
      n4059 <= 34'b0000000000000000000000000000000000;
    else
      n4059 <= n3300;
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:57:5  */
  assign n4060 = {n3333, port_out};
  /* ../../ext/neorv32/rtl/core/neorv32_gpio.vhd:140:5  */
  always @(posedge clk_i or posedge n3980)
    if (n3980)
      n4061 <= 1'b0;
    else
      n4061 <= n4038;
endmodule

module neorv32_boot_rom
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] );
  wire [79:0] n3190;
  wire [31:0] n3192;
  wire n3193;
  wire n3194;
  wire rden;
  wire [31:0] rdata;
  wire [4:0] n3197;
  wire [2:0] n3199;
  wire n3208;
  wire n3210;
  wire n3211;
  wire n3212;
  wire n3213;
  wire [31:0] n3218;
  reg n3221;
  wire [33:0] n3223;
  reg [31:0] n3227; // mem_rd
  assign \bus_rsp_o_bus_rsp_o[data]  = n3192; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n3193; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n3194; //(module output)
  assign n3190 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n3192 = n3223[31:0]; // extract
  assign n3193 = n3223[32]; // extract
  assign n3194 = n3223[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:38:10  */
  assign rden = n3221; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:39:10  */
  assign rdata = n3227; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:48:60  */
  assign n3197 = n3190[6:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:48:26  */
  assign n3199 = n3197[2:0];  // trunc
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:57:16  */
  assign n3208 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:60:25  */
  assign n3210 = n3190[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:60:48  */
  assign n3211 = n3190[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:60:34  */
  assign n3212 = ~n3211;
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:60:29  */
  assign n3213 = n3210 & n3212;
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:64:27  */
  assign n3218 = rden ? rdata : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:59:5  */
  always @(posedge clk_i or posedge n3208)
    if (n3208)
      n3221 <= 1'b0;
    else
      n3221 <= n3213;
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:47:5  */
  assign n3223 = {1'b0, rden, n3218};
  /* ../../ext/neorv32/rtl/core/neorv32_boot_rom.vhd:48:26  */
  reg [31:0] n3224[7:0] ; // memory
  initial begin
    n3224[7] = 32'b00000000000000000000000000000000;
    n3224[6] = 32'b00000000000000000000000000000000;
    n3224[5] = 32'b00000000000000101000000001100111;
    n3224[4] = 32'b11100000000000000000001010110111;
    n3224[3] = 32'b00000000111101110010000000100011;
    n3224[2] = 32'b01100000000101111000011110010011;
    n3224[1] = 32'b11111111111011110000011100110111;
    n3224[0] = 32'b00000000001000000111011110110111;
    end
  always @(posedge clk_i)
    if (1'b1)
      n3227 <= n3224[n3199];
endmodule

module neorv32_bus_io_switch_65536_19a0518872770ca4a65ad41d181dd3070f957778
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \main_req_i_main_req_i[addr] ,
   input  [31:0] \main_req_i_main_req_i[data] ,
   input  [3:0] \main_req_i_main_req_i[ben] ,
   input  \main_req_i_main_req_i[stb] ,
   input  \main_req_i_main_req_i[rw] ,
   input  \main_req_i_main_req_i[src] ,
   input  \main_req_i_main_req_i[priv] ,
   input  \main_req_i_main_req_i[amo] ,
   input  [3:0] \main_req_i_main_req_i[amoop] ,
   input  \main_req_i_main_req_i[fence] ,
   input  \main_req_i_main_req_i[sleep] ,
   input  \main_req_i_main_req_i[debug] ,
   input  [31:0] \dev_00_rsp_i_dev_00_rsp_i[data] ,
   input  \dev_00_rsp_i_dev_00_rsp_i[ack] ,
   input  \dev_00_rsp_i_dev_00_rsp_i[err] ,
   input  [31:0] \dev_01_rsp_i_dev_01_rsp_i[data] ,
   input  \dev_01_rsp_i_dev_01_rsp_i[ack] ,
   input  \dev_01_rsp_i_dev_01_rsp_i[err] ,
   input  [31:0] \dev_02_rsp_i_dev_02_rsp_i[data] ,
   input  \dev_02_rsp_i_dev_02_rsp_i[ack] ,
   input  \dev_02_rsp_i_dev_02_rsp_i[err] ,
   input  [31:0] \dev_03_rsp_i_dev_03_rsp_i[data] ,
   input  \dev_03_rsp_i_dev_03_rsp_i[ack] ,
   input  \dev_03_rsp_i_dev_03_rsp_i[err] ,
   input  [31:0] \dev_04_rsp_i_dev_04_rsp_i[data] ,
   input  \dev_04_rsp_i_dev_04_rsp_i[ack] ,
   input  \dev_04_rsp_i_dev_04_rsp_i[err] ,
   input  [31:0] \dev_05_rsp_i_dev_05_rsp_i[data] ,
   input  \dev_05_rsp_i_dev_05_rsp_i[ack] ,
   input  \dev_05_rsp_i_dev_05_rsp_i[err] ,
   input  [31:0] \dev_06_rsp_i_dev_06_rsp_i[data] ,
   input  \dev_06_rsp_i_dev_06_rsp_i[ack] ,
   input  \dev_06_rsp_i_dev_06_rsp_i[err] ,
   input  [31:0] \dev_07_rsp_i_dev_07_rsp_i[data] ,
   input  \dev_07_rsp_i_dev_07_rsp_i[ack] ,
   input  \dev_07_rsp_i_dev_07_rsp_i[err] ,
   input  [31:0] \dev_08_rsp_i_dev_08_rsp_i[data] ,
   input  \dev_08_rsp_i_dev_08_rsp_i[ack] ,
   input  \dev_08_rsp_i_dev_08_rsp_i[err] ,
   input  [31:0] \dev_09_rsp_i_dev_09_rsp_i[data] ,
   input  \dev_09_rsp_i_dev_09_rsp_i[ack] ,
   input  \dev_09_rsp_i_dev_09_rsp_i[err] ,
   input  [31:0] \dev_10_rsp_i_dev_10_rsp_i[data] ,
   input  \dev_10_rsp_i_dev_10_rsp_i[ack] ,
   input  \dev_10_rsp_i_dev_10_rsp_i[err] ,
   input  [31:0] \dev_11_rsp_i_dev_11_rsp_i[data] ,
   input  \dev_11_rsp_i_dev_11_rsp_i[ack] ,
   input  \dev_11_rsp_i_dev_11_rsp_i[err] ,
   input  [31:0] \dev_12_rsp_i_dev_12_rsp_i[data] ,
   input  \dev_12_rsp_i_dev_12_rsp_i[ack] ,
   input  \dev_12_rsp_i_dev_12_rsp_i[err] ,
   input  [31:0] \dev_13_rsp_i_dev_13_rsp_i[data] ,
   input  \dev_13_rsp_i_dev_13_rsp_i[ack] ,
   input  \dev_13_rsp_i_dev_13_rsp_i[err] ,
   input  [31:0] \dev_14_rsp_i_dev_14_rsp_i[data] ,
   input  \dev_14_rsp_i_dev_14_rsp_i[ack] ,
   input  \dev_14_rsp_i_dev_14_rsp_i[err] ,
   input  [31:0] \dev_15_rsp_i_dev_15_rsp_i[data] ,
   input  \dev_15_rsp_i_dev_15_rsp_i[ack] ,
   input  \dev_15_rsp_i_dev_15_rsp_i[err] ,
   input  [31:0] \dev_16_rsp_i_dev_16_rsp_i[data] ,
   input  \dev_16_rsp_i_dev_16_rsp_i[ack] ,
   input  \dev_16_rsp_i_dev_16_rsp_i[err] ,
   input  [31:0] \dev_17_rsp_i_dev_17_rsp_i[data] ,
   input  \dev_17_rsp_i_dev_17_rsp_i[ack] ,
   input  \dev_17_rsp_i_dev_17_rsp_i[err] ,
   input  [31:0] \dev_18_rsp_i_dev_18_rsp_i[data] ,
   input  \dev_18_rsp_i_dev_18_rsp_i[ack] ,
   input  \dev_18_rsp_i_dev_18_rsp_i[err] ,
   input  [31:0] \dev_19_rsp_i_dev_19_rsp_i[data] ,
   input  \dev_19_rsp_i_dev_19_rsp_i[ack] ,
   input  \dev_19_rsp_i_dev_19_rsp_i[err] ,
   input  [31:0] \dev_20_rsp_i_dev_20_rsp_i[data] ,
   input  \dev_20_rsp_i_dev_20_rsp_i[ack] ,
   input  \dev_20_rsp_i_dev_20_rsp_i[err] ,
   input  [31:0] \dev_21_rsp_i_dev_21_rsp_i[data] ,
   input  \dev_21_rsp_i_dev_21_rsp_i[ack] ,
   input  \dev_21_rsp_i_dev_21_rsp_i[err] ,
   input  [31:0] \dev_22_rsp_i_dev_22_rsp_i[data] ,
   input  \dev_22_rsp_i_dev_22_rsp_i[ack] ,
   input  \dev_22_rsp_i_dev_22_rsp_i[err] ,
   input  [31:0] \dev_23_rsp_i_dev_23_rsp_i[data] ,
   input  \dev_23_rsp_i_dev_23_rsp_i[ack] ,
   input  \dev_23_rsp_i_dev_23_rsp_i[err] ,
   input  [31:0] \dev_24_rsp_i_dev_24_rsp_i[data] ,
   input  \dev_24_rsp_i_dev_24_rsp_i[ack] ,
   input  \dev_24_rsp_i_dev_24_rsp_i[err] ,
   input  [31:0] \dev_25_rsp_i_dev_25_rsp_i[data] ,
   input  \dev_25_rsp_i_dev_25_rsp_i[ack] ,
   input  \dev_25_rsp_i_dev_25_rsp_i[err] ,
   input  [31:0] \dev_26_rsp_i_dev_26_rsp_i[data] ,
   input  \dev_26_rsp_i_dev_26_rsp_i[ack] ,
   input  \dev_26_rsp_i_dev_26_rsp_i[err] ,
   input  [31:0] \dev_27_rsp_i_dev_27_rsp_i[data] ,
   input  \dev_27_rsp_i_dev_27_rsp_i[ack] ,
   input  \dev_27_rsp_i_dev_27_rsp_i[err] ,
   input  [31:0] \dev_28_rsp_i_dev_28_rsp_i[data] ,
   input  \dev_28_rsp_i_dev_28_rsp_i[ack] ,
   input  \dev_28_rsp_i_dev_28_rsp_i[err] ,
   input  [31:0] \dev_29_rsp_i_dev_29_rsp_i[data] ,
   input  \dev_29_rsp_i_dev_29_rsp_i[ack] ,
   input  \dev_29_rsp_i_dev_29_rsp_i[err] ,
   input  [31:0] \dev_30_rsp_i_dev_30_rsp_i[data] ,
   input  \dev_30_rsp_i_dev_30_rsp_i[ack] ,
   input  \dev_30_rsp_i_dev_30_rsp_i[err] ,
   input  [31:0] \dev_31_rsp_i_dev_31_rsp_i[data] ,
   input  \dev_31_rsp_i_dev_31_rsp_i[ack] ,
   input  \dev_31_rsp_i_dev_31_rsp_i[err] ,
   output [31:0] \main_rsp_o_main_rsp_o[data] ,
   output \main_rsp_o_main_rsp_o[ack] ,
   output \main_rsp_o_main_rsp_o[err] ,
   output [31:0] \dev_00_req_o_dev_00_req_o[addr] ,
   output [31:0] \dev_00_req_o_dev_00_req_o[data] ,
   output [3:0] \dev_00_req_o_dev_00_req_o[ben] ,
   output \dev_00_req_o_dev_00_req_o[stb] ,
   output \dev_00_req_o_dev_00_req_o[rw] ,
   output \dev_00_req_o_dev_00_req_o[src] ,
   output \dev_00_req_o_dev_00_req_o[priv] ,
   output \dev_00_req_o_dev_00_req_o[amo] ,
   output [3:0] \dev_00_req_o_dev_00_req_o[amoop] ,
   output \dev_00_req_o_dev_00_req_o[fence] ,
   output \dev_00_req_o_dev_00_req_o[sleep] ,
   output \dev_00_req_o_dev_00_req_o[debug] ,
   output [31:0] \dev_01_req_o_dev_01_req_o[addr] ,
   output [31:0] \dev_01_req_o_dev_01_req_o[data] ,
   output [3:0] \dev_01_req_o_dev_01_req_o[ben] ,
   output \dev_01_req_o_dev_01_req_o[stb] ,
   output \dev_01_req_o_dev_01_req_o[rw] ,
   output \dev_01_req_o_dev_01_req_o[src] ,
   output \dev_01_req_o_dev_01_req_o[priv] ,
   output \dev_01_req_o_dev_01_req_o[amo] ,
   output [3:0] \dev_01_req_o_dev_01_req_o[amoop] ,
   output \dev_01_req_o_dev_01_req_o[fence] ,
   output \dev_01_req_o_dev_01_req_o[sleep] ,
   output \dev_01_req_o_dev_01_req_o[debug] ,
   output [31:0] \dev_02_req_o_dev_02_req_o[addr] ,
   output [31:0] \dev_02_req_o_dev_02_req_o[data] ,
   output [3:0] \dev_02_req_o_dev_02_req_o[ben] ,
   output \dev_02_req_o_dev_02_req_o[stb] ,
   output \dev_02_req_o_dev_02_req_o[rw] ,
   output \dev_02_req_o_dev_02_req_o[src] ,
   output \dev_02_req_o_dev_02_req_o[priv] ,
   output \dev_02_req_o_dev_02_req_o[amo] ,
   output [3:0] \dev_02_req_o_dev_02_req_o[amoop] ,
   output \dev_02_req_o_dev_02_req_o[fence] ,
   output \dev_02_req_o_dev_02_req_o[sleep] ,
   output \dev_02_req_o_dev_02_req_o[debug] ,
   output [31:0] \dev_03_req_o_dev_03_req_o[addr] ,
   output [31:0] \dev_03_req_o_dev_03_req_o[data] ,
   output [3:0] \dev_03_req_o_dev_03_req_o[ben] ,
   output \dev_03_req_o_dev_03_req_o[stb] ,
   output \dev_03_req_o_dev_03_req_o[rw] ,
   output \dev_03_req_o_dev_03_req_o[src] ,
   output \dev_03_req_o_dev_03_req_o[priv] ,
   output \dev_03_req_o_dev_03_req_o[amo] ,
   output [3:0] \dev_03_req_o_dev_03_req_o[amoop] ,
   output \dev_03_req_o_dev_03_req_o[fence] ,
   output \dev_03_req_o_dev_03_req_o[sleep] ,
   output \dev_03_req_o_dev_03_req_o[debug] ,
   output [31:0] \dev_04_req_o_dev_04_req_o[addr] ,
   output [31:0] \dev_04_req_o_dev_04_req_o[data] ,
   output [3:0] \dev_04_req_o_dev_04_req_o[ben] ,
   output \dev_04_req_o_dev_04_req_o[stb] ,
   output \dev_04_req_o_dev_04_req_o[rw] ,
   output \dev_04_req_o_dev_04_req_o[src] ,
   output \dev_04_req_o_dev_04_req_o[priv] ,
   output \dev_04_req_o_dev_04_req_o[amo] ,
   output [3:0] \dev_04_req_o_dev_04_req_o[amoop] ,
   output \dev_04_req_o_dev_04_req_o[fence] ,
   output \dev_04_req_o_dev_04_req_o[sleep] ,
   output \dev_04_req_o_dev_04_req_o[debug] ,
   output [31:0] \dev_05_req_o_dev_05_req_o[addr] ,
   output [31:0] \dev_05_req_o_dev_05_req_o[data] ,
   output [3:0] \dev_05_req_o_dev_05_req_o[ben] ,
   output \dev_05_req_o_dev_05_req_o[stb] ,
   output \dev_05_req_o_dev_05_req_o[rw] ,
   output \dev_05_req_o_dev_05_req_o[src] ,
   output \dev_05_req_o_dev_05_req_o[priv] ,
   output \dev_05_req_o_dev_05_req_o[amo] ,
   output [3:0] \dev_05_req_o_dev_05_req_o[amoop] ,
   output \dev_05_req_o_dev_05_req_o[fence] ,
   output \dev_05_req_o_dev_05_req_o[sleep] ,
   output \dev_05_req_o_dev_05_req_o[debug] ,
   output [31:0] \dev_06_req_o_dev_06_req_o[addr] ,
   output [31:0] \dev_06_req_o_dev_06_req_o[data] ,
   output [3:0] \dev_06_req_o_dev_06_req_o[ben] ,
   output \dev_06_req_o_dev_06_req_o[stb] ,
   output \dev_06_req_o_dev_06_req_o[rw] ,
   output \dev_06_req_o_dev_06_req_o[src] ,
   output \dev_06_req_o_dev_06_req_o[priv] ,
   output \dev_06_req_o_dev_06_req_o[amo] ,
   output [3:0] \dev_06_req_o_dev_06_req_o[amoop] ,
   output \dev_06_req_o_dev_06_req_o[fence] ,
   output \dev_06_req_o_dev_06_req_o[sleep] ,
   output \dev_06_req_o_dev_06_req_o[debug] ,
   output [31:0] \dev_07_req_o_dev_07_req_o[addr] ,
   output [31:0] \dev_07_req_o_dev_07_req_o[data] ,
   output [3:0] \dev_07_req_o_dev_07_req_o[ben] ,
   output \dev_07_req_o_dev_07_req_o[stb] ,
   output \dev_07_req_o_dev_07_req_o[rw] ,
   output \dev_07_req_o_dev_07_req_o[src] ,
   output \dev_07_req_o_dev_07_req_o[priv] ,
   output \dev_07_req_o_dev_07_req_o[amo] ,
   output [3:0] \dev_07_req_o_dev_07_req_o[amoop] ,
   output \dev_07_req_o_dev_07_req_o[fence] ,
   output \dev_07_req_o_dev_07_req_o[sleep] ,
   output \dev_07_req_o_dev_07_req_o[debug] ,
   output [31:0] \dev_08_req_o_dev_08_req_o[addr] ,
   output [31:0] \dev_08_req_o_dev_08_req_o[data] ,
   output [3:0] \dev_08_req_o_dev_08_req_o[ben] ,
   output \dev_08_req_o_dev_08_req_o[stb] ,
   output \dev_08_req_o_dev_08_req_o[rw] ,
   output \dev_08_req_o_dev_08_req_o[src] ,
   output \dev_08_req_o_dev_08_req_o[priv] ,
   output \dev_08_req_o_dev_08_req_o[amo] ,
   output [3:0] \dev_08_req_o_dev_08_req_o[amoop] ,
   output \dev_08_req_o_dev_08_req_o[fence] ,
   output \dev_08_req_o_dev_08_req_o[sleep] ,
   output \dev_08_req_o_dev_08_req_o[debug] ,
   output [31:0] \dev_09_req_o_dev_09_req_o[addr] ,
   output [31:0] \dev_09_req_o_dev_09_req_o[data] ,
   output [3:0] \dev_09_req_o_dev_09_req_o[ben] ,
   output \dev_09_req_o_dev_09_req_o[stb] ,
   output \dev_09_req_o_dev_09_req_o[rw] ,
   output \dev_09_req_o_dev_09_req_o[src] ,
   output \dev_09_req_o_dev_09_req_o[priv] ,
   output \dev_09_req_o_dev_09_req_o[amo] ,
   output [3:0] \dev_09_req_o_dev_09_req_o[amoop] ,
   output \dev_09_req_o_dev_09_req_o[fence] ,
   output \dev_09_req_o_dev_09_req_o[sleep] ,
   output \dev_09_req_o_dev_09_req_o[debug] ,
   output [31:0] \dev_10_req_o_dev_10_req_o[addr] ,
   output [31:0] \dev_10_req_o_dev_10_req_o[data] ,
   output [3:0] \dev_10_req_o_dev_10_req_o[ben] ,
   output \dev_10_req_o_dev_10_req_o[stb] ,
   output \dev_10_req_o_dev_10_req_o[rw] ,
   output \dev_10_req_o_dev_10_req_o[src] ,
   output \dev_10_req_o_dev_10_req_o[priv] ,
   output \dev_10_req_o_dev_10_req_o[amo] ,
   output [3:0] \dev_10_req_o_dev_10_req_o[amoop] ,
   output \dev_10_req_o_dev_10_req_o[fence] ,
   output \dev_10_req_o_dev_10_req_o[sleep] ,
   output \dev_10_req_o_dev_10_req_o[debug] ,
   output [31:0] \dev_11_req_o_dev_11_req_o[addr] ,
   output [31:0] \dev_11_req_o_dev_11_req_o[data] ,
   output [3:0] \dev_11_req_o_dev_11_req_o[ben] ,
   output \dev_11_req_o_dev_11_req_o[stb] ,
   output \dev_11_req_o_dev_11_req_o[rw] ,
   output \dev_11_req_o_dev_11_req_o[src] ,
   output \dev_11_req_o_dev_11_req_o[priv] ,
   output \dev_11_req_o_dev_11_req_o[amo] ,
   output [3:0] \dev_11_req_o_dev_11_req_o[amoop] ,
   output \dev_11_req_o_dev_11_req_o[fence] ,
   output \dev_11_req_o_dev_11_req_o[sleep] ,
   output \dev_11_req_o_dev_11_req_o[debug] ,
   output [31:0] \dev_12_req_o_dev_12_req_o[addr] ,
   output [31:0] \dev_12_req_o_dev_12_req_o[data] ,
   output [3:0] \dev_12_req_o_dev_12_req_o[ben] ,
   output \dev_12_req_o_dev_12_req_o[stb] ,
   output \dev_12_req_o_dev_12_req_o[rw] ,
   output \dev_12_req_o_dev_12_req_o[src] ,
   output \dev_12_req_o_dev_12_req_o[priv] ,
   output \dev_12_req_o_dev_12_req_o[amo] ,
   output [3:0] \dev_12_req_o_dev_12_req_o[amoop] ,
   output \dev_12_req_o_dev_12_req_o[fence] ,
   output \dev_12_req_o_dev_12_req_o[sleep] ,
   output \dev_12_req_o_dev_12_req_o[debug] ,
   output [31:0] \dev_13_req_o_dev_13_req_o[addr] ,
   output [31:0] \dev_13_req_o_dev_13_req_o[data] ,
   output [3:0] \dev_13_req_o_dev_13_req_o[ben] ,
   output \dev_13_req_o_dev_13_req_o[stb] ,
   output \dev_13_req_o_dev_13_req_o[rw] ,
   output \dev_13_req_o_dev_13_req_o[src] ,
   output \dev_13_req_o_dev_13_req_o[priv] ,
   output \dev_13_req_o_dev_13_req_o[amo] ,
   output [3:0] \dev_13_req_o_dev_13_req_o[amoop] ,
   output \dev_13_req_o_dev_13_req_o[fence] ,
   output \dev_13_req_o_dev_13_req_o[sleep] ,
   output \dev_13_req_o_dev_13_req_o[debug] ,
   output [31:0] \dev_14_req_o_dev_14_req_o[addr] ,
   output [31:0] \dev_14_req_o_dev_14_req_o[data] ,
   output [3:0] \dev_14_req_o_dev_14_req_o[ben] ,
   output \dev_14_req_o_dev_14_req_o[stb] ,
   output \dev_14_req_o_dev_14_req_o[rw] ,
   output \dev_14_req_o_dev_14_req_o[src] ,
   output \dev_14_req_o_dev_14_req_o[priv] ,
   output \dev_14_req_o_dev_14_req_o[amo] ,
   output [3:0] \dev_14_req_o_dev_14_req_o[amoop] ,
   output \dev_14_req_o_dev_14_req_o[fence] ,
   output \dev_14_req_o_dev_14_req_o[sleep] ,
   output \dev_14_req_o_dev_14_req_o[debug] ,
   output [31:0] \dev_15_req_o_dev_15_req_o[addr] ,
   output [31:0] \dev_15_req_o_dev_15_req_o[data] ,
   output [3:0] \dev_15_req_o_dev_15_req_o[ben] ,
   output \dev_15_req_o_dev_15_req_o[stb] ,
   output \dev_15_req_o_dev_15_req_o[rw] ,
   output \dev_15_req_o_dev_15_req_o[src] ,
   output \dev_15_req_o_dev_15_req_o[priv] ,
   output \dev_15_req_o_dev_15_req_o[amo] ,
   output [3:0] \dev_15_req_o_dev_15_req_o[amoop] ,
   output \dev_15_req_o_dev_15_req_o[fence] ,
   output \dev_15_req_o_dev_15_req_o[sleep] ,
   output \dev_15_req_o_dev_15_req_o[debug] ,
   output [31:0] \dev_16_req_o_dev_16_req_o[addr] ,
   output [31:0] \dev_16_req_o_dev_16_req_o[data] ,
   output [3:0] \dev_16_req_o_dev_16_req_o[ben] ,
   output \dev_16_req_o_dev_16_req_o[stb] ,
   output \dev_16_req_o_dev_16_req_o[rw] ,
   output \dev_16_req_o_dev_16_req_o[src] ,
   output \dev_16_req_o_dev_16_req_o[priv] ,
   output \dev_16_req_o_dev_16_req_o[amo] ,
   output [3:0] \dev_16_req_o_dev_16_req_o[amoop] ,
   output \dev_16_req_o_dev_16_req_o[fence] ,
   output \dev_16_req_o_dev_16_req_o[sleep] ,
   output \dev_16_req_o_dev_16_req_o[debug] ,
   output [31:0] \dev_17_req_o_dev_17_req_o[addr] ,
   output [31:0] \dev_17_req_o_dev_17_req_o[data] ,
   output [3:0] \dev_17_req_o_dev_17_req_o[ben] ,
   output \dev_17_req_o_dev_17_req_o[stb] ,
   output \dev_17_req_o_dev_17_req_o[rw] ,
   output \dev_17_req_o_dev_17_req_o[src] ,
   output \dev_17_req_o_dev_17_req_o[priv] ,
   output \dev_17_req_o_dev_17_req_o[amo] ,
   output [3:0] \dev_17_req_o_dev_17_req_o[amoop] ,
   output \dev_17_req_o_dev_17_req_o[fence] ,
   output \dev_17_req_o_dev_17_req_o[sleep] ,
   output \dev_17_req_o_dev_17_req_o[debug] ,
   output [31:0] \dev_18_req_o_dev_18_req_o[addr] ,
   output [31:0] \dev_18_req_o_dev_18_req_o[data] ,
   output [3:0] \dev_18_req_o_dev_18_req_o[ben] ,
   output \dev_18_req_o_dev_18_req_o[stb] ,
   output \dev_18_req_o_dev_18_req_o[rw] ,
   output \dev_18_req_o_dev_18_req_o[src] ,
   output \dev_18_req_o_dev_18_req_o[priv] ,
   output \dev_18_req_o_dev_18_req_o[amo] ,
   output [3:0] \dev_18_req_o_dev_18_req_o[amoop] ,
   output \dev_18_req_o_dev_18_req_o[fence] ,
   output \dev_18_req_o_dev_18_req_o[sleep] ,
   output \dev_18_req_o_dev_18_req_o[debug] ,
   output [31:0] \dev_19_req_o_dev_19_req_o[addr] ,
   output [31:0] \dev_19_req_o_dev_19_req_o[data] ,
   output [3:0] \dev_19_req_o_dev_19_req_o[ben] ,
   output \dev_19_req_o_dev_19_req_o[stb] ,
   output \dev_19_req_o_dev_19_req_o[rw] ,
   output \dev_19_req_o_dev_19_req_o[src] ,
   output \dev_19_req_o_dev_19_req_o[priv] ,
   output \dev_19_req_o_dev_19_req_o[amo] ,
   output [3:0] \dev_19_req_o_dev_19_req_o[amoop] ,
   output \dev_19_req_o_dev_19_req_o[fence] ,
   output \dev_19_req_o_dev_19_req_o[sleep] ,
   output \dev_19_req_o_dev_19_req_o[debug] ,
   output [31:0] \dev_20_req_o_dev_20_req_o[addr] ,
   output [31:0] \dev_20_req_o_dev_20_req_o[data] ,
   output [3:0] \dev_20_req_o_dev_20_req_o[ben] ,
   output \dev_20_req_o_dev_20_req_o[stb] ,
   output \dev_20_req_o_dev_20_req_o[rw] ,
   output \dev_20_req_o_dev_20_req_o[src] ,
   output \dev_20_req_o_dev_20_req_o[priv] ,
   output \dev_20_req_o_dev_20_req_o[amo] ,
   output [3:0] \dev_20_req_o_dev_20_req_o[amoop] ,
   output \dev_20_req_o_dev_20_req_o[fence] ,
   output \dev_20_req_o_dev_20_req_o[sleep] ,
   output \dev_20_req_o_dev_20_req_o[debug] ,
   output [31:0] \dev_21_req_o_dev_21_req_o[addr] ,
   output [31:0] \dev_21_req_o_dev_21_req_o[data] ,
   output [3:0] \dev_21_req_o_dev_21_req_o[ben] ,
   output \dev_21_req_o_dev_21_req_o[stb] ,
   output \dev_21_req_o_dev_21_req_o[rw] ,
   output \dev_21_req_o_dev_21_req_o[src] ,
   output \dev_21_req_o_dev_21_req_o[priv] ,
   output \dev_21_req_o_dev_21_req_o[amo] ,
   output [3:0] \dev_21_req_o_dev_21_req_o[amoop] ,
   output \dev_21_req_o_dev_21_req_o[fence] ,
   output \dev_21_req_o_dev_21_req_o[sleep] ,
   output \dev_21_req_o_dev_21_req_o[debug] ,
   output [31:0] \dev_22_req_o_dev_22_req_o[addr] ,
   output [31:0] \dev_22_req_o_dev_22_req_o[data] ,
   output [3:0] \dev_22_req_o_dev_22_req_o[ben] ,
   output \dev_22_req_o_dev_22_req_o[stb] ,
   output \dev_22_req_o_dev_22_req_o[rw] ,
   output \dev_22_req_o_dev_22_req_o[src] ,
   output \dev_22_req_o_dev_22_req_o[priv] ,
   output \dev_22_req_o_dev_22_req_o[amo] ,
   output [3:0] \dev_22_req_o_dev_22_req_o[amoop] ,
   output \dev_22_req_o_dev_22_req_o[fence] ,
   output \dev_22_req_o_dev_22_req_o[sleep] ,
   output \dev_22_req_o_dev_22_req_o[debug] ,
   output [31:0] \dev_23_req_o_dev_23_req_o[addr] ,
   output [31:0] \dev_23_req_o_dev_23_req_o[data] ,
   output [3:0] \dev_23_req_o_dev_23_req_o[ben] ,
   output \dev_23_req_o_dev_23_req_o[stb] ,
   output \dev_23_req_o_dev_23_req_o[rw] ,
   output \dev_23_req_o_dev_23_req_o[src] ,
   output \dev_23_req_o_dev_23_req_o[priv] ,
   output \dev_23_req_o_dev_23_req_o[amo] ,
   output [3:0] \dev_23_req_o_dev_23_req_o[amoop] ,
   output \dev_23_req_o_dev_23_req_o[fence] ,
   output \dev_23_req_o_dev_23_req_o[sleep] ,
   output \dev_23_req_o_dev_23_req_o[debug] ,
   output [31:0] \dev_24_req_o_dev_24_req_o[addr] ,
   output [31:0] \dev_24_req_o_dev_24_req_o[data] ,
   output [3:0] \dev_24_req_o_dev_24_req_o[ben] ,
   output \dev_24_req_o_dev_24_req_o[stb] ,
   output \dev_24_req_o_dev_24_req_o[rw] ,
   output \dev_24_req_o_dev_24_req_o[src] ,
   output \dev_24_req_o_dev_24_req_o[priv] ,
   output \dev_24_req_o_dev_24_req_o[amo] ,
   output [3:0] \dev_24_req_o_dev_24_req_o[amoop] ,
   output \dev_24_req_o_dev_24_req_o[fence] ,
   output \dev_24_req_o_dev_24_req_o[sleep] ,
   output \dev_24_req_o_dev_24_req_o[debug] ,
   output [31:0] \dev_25_req_o_dev_25_req_o[addr] ,
   output [31:0] \dev_25_req_o_dev_25_req_o[data] ,
   output [3:0] \dev_25_req_o_dev_25_req_o[ben] ,
   output \dev_25_req_o_dev_25_req_o[stb] ,
   output \dev_25_req_o_dev_25_req_o[rw] ,
   output \dev_25_req_o_dev_25_req_o[src] ,
   output \dev_25_req_o_dev_25_req_o[priv] ,
   output \dev_25_req_o_dev_25_req_o[amo] ,
   output [3:0] \dev_25_req_o_dev_25_req_o[amoop] ,
   output \dev_25_req_o_dev_25_req_o[fence] ,
   output \dev_25_req_o_dev_25_req_o[sleep] ,
   output \dev_25_req_o_dev_25_req_o[debug] ,
   output [31:0] \dev_26_req_o_dev_26_req_o[addr] ,
   output [31:0] \dev_26_req_o_dev_26_req_o[data] ,
   output [3:0] \dev_26_req_o_dev_26_req_o[ben] ,
   output \dev_26_req_o_dev_26_req_o[stb] ,
   output \dev_26_req_o_dev_26_req_o[rw] ,
   output \dev_26_req_o_dev_26_req_o[src] ,
   output \dev_26_req_o_dev_26_req_o[priv] ,
   output \dev_26_req_o_dev_26_req_o[amo] ,
   output [3:0] \dev_26_req_o_dev_26_req_o[amoop] ,
   output \dev_26_req_o_dev_26_req_o[fence] ,
   output \dev_26_req_o_dev_26_req_o[sleep] ,
   output \dev_26_req_o_dev_26_req_o[debug] ,
   output [31:0] \dev_27_req_o_dev_27_req_o[addr] ,
   output [31:0] \dev_27_req_o_dev_27_req_o[data] ,
   output [3:0] \dev_27_req_o_dev_27_req_o[ben] ,
   output \dev_27_req_o_dev_27_req_o[stb] ,
   output \dev_27_req_o_dev_27_req_o[rw] ,
   output \dev_27_req_o_dev_27_req_o[src] ,
   output \dev_27_req_o_dev_27_req_o[priv] ,
   output \dev_27_req_o_dev_27_req_o[amo] ,
   output [3:0] \dev_27_req_o_dev_27_req_o[amoop] ,
   output \dev_27_req_o_dev_27_req_o[fence] ,
   output \dev_27_req_o_dev_27_req_o[sleep] ,
   output \dev_27_req_o_dev_27_req_o[debug] ,
   output [31:0] \dev_28_req_o_dev_28_req_o[addr] ,
   output [31:0] \dev_28_req_o_dev_28_req_o[data] ,
   output [3:0] \dev_28_req_o_dev_28_req_o[ben] ,
   output \dev_28_req_o_dev_28_req_o[stb] ,
   output \dev_28_req_o_dev_28_req_o[rw] ,
   output \dev_28_req_o_dev_28_req_o[src] ,
   output \dev_28_req_o_dev_28_req_o[priv] ,
   output \dev_28_req_o_dev_28_req_o[amo] ,
   output [3:0] \dev_28_req_o_dev_28_req_o[amoop] ,
   output \dev_28_req_o_dev_28_req_o[fence] ,
   output \dev_28_req_o_dev_28_req_o[sleep] ,
   output \dev_28_req_o_dev_28_req_o[debug] ,
   output [31:0] \dev_29_req_o_dev_29_req_o[addr] ,
   output [31:0] \dev_29_req_o_dev_29_req_o[data] ,
   output [3:0] \dev_29_req_o_dev_29_req_o[ben] ,
   output \dev_29_req_o_dev_29_req_o[stb] ,
   output \dev_29_req_o_dev_29_req_o[rw] ,
   output \dev_29_req_o_dev_29_req_o[src] ,
   output \dev_29_req_o_dev_29_req_o[priv] ,
   output \dev_29_req_o_dev_29_req_o[amo] ,
   output [3:0] \dev_29_req_o_dev_29_req_o[amoop] ,
   output \dev_29_req_o_dev_29_req_o[fence] ,
   output \dev_29_req_o_dev_29_req_o[sleep] ,
   output \dev_29_req_o_dev_29_req_o[debug] ,
   output [31:0] \dev_30_req_o_dev_30_req_o[addr] ,
   output [31:0] \dev_30_req_o_dev_30_req_o[data] ,
   output [3:0] \dev_30_req_o_dev_30_req_o[ben] ,
   output \dev_30_req_o_dev_30_req_o[stb] ,
   output \dev_30_req_o_dev_30_req_o[rw] ,
   output \dev_30_req_o_dev_30_req_o[src] ,
   output \dev_30_req_o_dev_30_req_o[priv] ,
   output \dev_30_req_o_dev_30_req_o[amo] ,
   output [3:0] \dev_30_req_o_dev_30_req_o[amoop] ,
   output \dev_30_req_o_dev_30_req_o[fence] ,
   output \dev_30_req_o_dev_30_req_o[sleep] ,
   output \dev_30_req_o_dev_30_req_o[debug] ,
   output [31:0] \dev_31_req_o_dev_31_req_o[addr] ,
   output [31:0] \dev_31_req_o_dev_31_req_o[data] ,
   output [3:0] \dev_31_req_o_dev_31_req_o[ben] ,
   output \dev_31_req_o_dev_31_req_o[stb] ,
   output \dev_31_req_o_dev_31_req_o[rw] ,
   output \dev_31_req_o_dev_31_req_o[src] ,
   output \dev_31_req_o_dev_31_req_o[priv] ,
   output \dev_31_req_o_dev_31_req_o[amo] ,
   output [3:0] \dev_31_req_o_dev_31_req_o[amoop] ,
   output \dev_31_req_o_dev_31_req_o[fence] ,
   output \dev_31_req_o_dev_31_req_o[sleep] ,
   output \dev_31_req_o_dev_31_req_o[debug] );
  wire [79:0] n2421;
  wire [31:0] n2423;
  wire n2424;
  wire n2425;
  wire [31:0] n2427;
  wire [31:0] n2428;
  wire [3:0] n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire [3:0] n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire [33:0] n2439;
  wire [31:0] n2441;
  wire [31:0] n2442;
  wire [3:0] n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire [3:0] n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire [33:0] n2453;
  wire [31:0] n2455;
  wire [31:0] n2456;
  wire [3:0] n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire [3:0] n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire [33:0] n2467;
  wire [31:0] n2469;
  wire [31:0] n2470;
  wire [3:0] n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire [3:0] n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire [33:0] n2481;
  wire [31:0] n2483;
  wire [31:0] n2484;
  wire [3:0] n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire [3:0] n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire [33:0] n2495;
  wire [31:0] n2497;
  wire [31:0] n2498;
  wire [3:0] n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire [3:0] n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire [33:0] n2509;
  wire [31:0] n2511;
  wire [31:0] n2512;
  wire [3:0] n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire [3:0] n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire [33:0] n2523;
  wire [31:0] n2525;
  wire [31:0] n2526;
  wire [3:0] n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire [3:0] n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire [33:0] n2537;
  wire [31:0] n2539;
  wire [31:0] n2540;
  wire [3:0] n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire [3:0] n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire [33:0] n2551;
  wire [31:0] n2553;
  wire [31:0] n2554;
  wire [3:0] n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire [3:0] n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire [33:0] n2565;
  wire [31:0] n2567;
  wire [31:0] n2568;
  wire [3:0] n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire [3:0] n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire [33:0] n2579;
  wire [31:0] n2581;
  wire [31:0] n2582;
  wire [3:0] n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire [3:0] n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire [33:0] n2593;
  wire [31:0] n2595;
  wire [31:0] n2596;
  wire [3:0] n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire [3:0] n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire [33:0] n2607;
  wire [31:0] n2609;
  wire [31:0] n2610;
  wire [3:0] n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire [3:0] n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire [33:0] n2621;
  wire [31:0] n2623;
  wire [31:0] n2624;
  wire [3:0] n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire [3:0] n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire [33:0] n2635;
  wire [31:0] n2637;
  wire [31:0] n2638;
  wire [3:0] n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire [3:0] n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire [33:0] n2649;
  wire [31:0] n2651;
  wire [31:0] n2652;
  wire [3:0] n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire [3:0] n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire [33:0] n2663;
  wire [31:0] n2665;
  wire [31:0] n2666;
  wire [3:0] n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire [3:0] n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire [33:0] n2677;
  wire [31:0] n2679;
  wire [31:0] n2680;
  wire [3:0] n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire [3:0] n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire [33:0] n2691;
  wire [31:0] n2693;
  wire [31:0] n2694;
  wire [3:0] n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire [3:0] n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire [33:0] n2705;
  wire [31:0] n2707;
  wire [31:0] n2708;
  wire [3:0] n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire [3:0] n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire [33:0] n2719;
  wire [31:0] n2721;
  wire [31:0] n2722;
  wire [3:0] n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire [3:0] n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire [33:0] n2733;
  wire [31:0] n2735;
  wire [31:0] n2736;
  wire [3:0] n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire [3:0] n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire [33:0] n2747;
  wire [31:0] n2749;
  wire [31:0] n2750;
  wire [3:0] n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire [3:0] n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire [33:0] n2761;
  wire [31:0] n2763;
  wire [31:0] n2764;
  wire [3:0] n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire [3:0] n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire [33:0] n2775;
  wire [31:0] n2777;
  wire [31:0] n2778;
  wire [3:0] n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire [3:0] n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire [33:0] n2789;
  wire [31:0] n2791;
  wire [31:0] n2792;
  wire [3:0] n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire [3:0] n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire [33:0] n2803;
  wire [31:0] n2805;
  wire [31:0] n2806;
  wire [3:0] n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire [3:0] n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire [33:0] n2817;
  wire [31:0] n2819;
  wire [31:0] n2820;
  wire [3:0] n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire [3:0] n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire [33:0] n2831;
  wire [31:0] n2833;
  wire [31:0] n2834;
  wire [3:0] n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire [3:0] n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire [33:0] n2845;
  wire [31:0] n2847;
  wire [31:0] n2848;
  wire [3:0] n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire [3:0] n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire [33:0] n2859;
  wire [31:0] n2861;
  wire [31:0] n2862;
  wire [3:0] n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire [3:0] n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire [33:0] n2873;
  wire [2559:0] dev_req;
  wire [1087:0] dev_rsp;
  wire [79:0] main_req;
  wire [33:0] main_rsp;
  wire [33:0] neorv32_bus_reg_inst_n2874;
  wire [79:0] neorv32_bus_reg_inst_n2875;
  wire [31:0] \neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[data] ;
  wire \neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[ack] ;
  wire \neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[err] ;
  wire [31:0] \neorv32_bus_reg_inst.device_req_o_device_req_o[addr] ;
  wire [31:0] \neorv32_bus_reg_inst.device_req_o_device_req_o[data] ;
  wire [3:0] \neorv32_bus_reg_inst.device_req_o_device_req_o[ben] ;
  wire \neorv32_bus_reg_inst.device_req_o_device_req_o[stb] ;
  wire \neorv32_bus_reg_inst.device_req_o_device_req_o[rw] ;
  wire \neorv32_bus_reg_inst.device_req_o_device_req_o[src] ;
  wire \neorv32_bus_reg_inst.device_req_o_device_req_o[priv] ;
  wire \neorv32_bus_reg_inst.device_req_o_device_req_o[amo] ;
  wire [3:0] \neorv32_bus_reg_inst.device_req_o_device_req_o[amoop] ;
  wire \neorv32_bus_reg_inst.device_req_o_device_req_o[fence] ;
  wire \neorv32_bus_reg_inst.device_req_o_device_req_o[sleep] ;
  wire \neorv32_bus_reg_inst.device_req_o_device_req_o[debug] ;
  wire [31:0] n2876;
  wire [31:0] n2877;
  wire [3:0] n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire [3:0] n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire [33:0] n2888;
  wire [79:0] n2890;
  wire [31:0] n2892;
  wire n2893;
  wire n2894;
  wire [79:0] n2897;
  wire [79:0] n2898;
  wire [79:0] n2899;
  wire [79:0] n2900;
  wire [79:0] n2901;
  wire [79:0] n2902;
  wire [79:0] n2903;
  wire [79:0] n2904;
  wire [79:0] n2905;
  wire [79:0] n2906;
  wire [79:0] n2907;
  wire [79:0] n2908;
  wire [79:0] n2909;
  wire [79:0] n2910;
  wire [79:0] n2911;
  wire [79:0] n2912;
  wire [79:0] n2913;
  wire [79:0] n2914;
  wire [79:0] n2915;
  wire [79:0] n2916;
  wire [79:0] n2917;
  wire [79:0] n2918;
  wire [79:0] n2919;
  wire [79:0] n2920;
  wire [79:0] n2921;
  wire [79:0] n2922;
  wire [79:0] n2923;
  wire [79:0] n2924;
  wire [79:0] n2925;
  wire [79:0] n2926;
  wire [79:0] n2927;
  wire [79:0] n2928;
  wire [4:0] n2930;
  wire n2932;
  wire n2933;
  wire n2935;
  wire [10:0] n2936;
  wire [67:0] n2937;
  wire [4:0] n2941;
  wire n2943;
  wire n2944;
  wire n2946;
  wire [10:0] n2947;
  wire [67:0] n2948;
  wire [4:0] n2951;
  wire n2953;
  wire n2954;
  wire n2956;
  wire [10:0] n2957;
  wire [67:0] n2958;
  wire [4:0] n2961;
  wire n2963;
  wire n2964;
  wire n2966;
  wire [10:0] n2967;
  wire [67:0] n2968;
  wire [4:0] n2971;
  wire n2973;
  wire n2974;
  wire n2976;
  wire [10:0] n2977;
  wire [67:0] n2978;
  wire [4:0] n2981;
  wire n2983;
  wire n2984;
  wire n2986;
  wire [10:0] n2987;
  wire [67:0] n2988;
  wire [4:0] n2991;
  wire n2993;
  wire n2994;
  wire n2996;
  wire [10:0] n2997;
  wire [67:0] n2998;
  wire [4:0] n3001;
  wire n3003;
  wire n3004;
  wire n3006;
  wire [10:0] n3007;
  wire [67:0] n3008;
  wire [4:0] n3011;
  wire n3013;
  wire n3014;
  wire n3016;
  wire [10:0] n3017;
  wire [67:0] n3018;
  wire [4:0] n3021;
  wire n3023;
  wire n3024;
  wire n3026;
  wire [10:0] n3027;
  wire [67:0] n3028;
  localparam [33:0] n3032 = 34'b0000000000000000000000000000000000;
  wire [31:0] n3033;
  wire [31:0] n3035;
  wire [31:0] n3036;
  localparam [33:0] n3037 = 34'b0000000000000000000000000000000000;
  wire [1:0] n3038;
  wire [33:0] n3039;
  wire n3040;
  wire n3042;
  wire n3043;
  wire n3044;
  wire [33:0] n3045;
  wire n3046;
  wire n3048;
  wire n3049;
  wire [33:0] n3050;
  wire [31:0] n3051;
  wire [31:0] n3053;
  wire [31:0] n3054;
  wire [33:0] n3055;
  wire n3056;
  wire n3058;
  wire n3059;
  wire [33:0] n3060;
  wire n3061;
  wire n3063;
  wire n3064;
  wire [33:0] n3065;
  wire [31:0] n3066;
  wire [31:0] n3068;
  wire [31:0] n3069;
  wire [33:0] n3070;
  wire n3071;
  wire n3073;
  wire n3074;
  wire [33:0] n3075;
  wire n3076;
  wire n3078;
  wire n3079;
  wire [33:0] n3080;
  wire [31:0] n3081;
  wire [31:0] n3083;
  wire [31:0] n3084;
  wire [33:0] n3085;
  wire n3086;
  wire n3088;
  wire n3089;
  wire [33:0] n3090;
  wire n3091;
  wire n3093;
  wire n3094;
  wire [33:0] n3095;
  wire [31:0] n3096;
  wire [31:0] n3098;
  wire [31:0] n3099;
  wire [33:0] n3100;
  wire n3101;
  wire n3103;
  wire n3104;
  wire [33:0] n3105;
  wire n3106;
  wire n3108;
  wire n3109;
  wire [33:0] n3110;
  wire [31:0] n3111;
  wire [31:0] n3113;
  wire [31:0] n3114;
  wire [33:0] n3115;
  wire n3116;
  wire n3118;
  wire n3119;
  wire [33:0] n3120;
  wire n3121;
  wire n3123;
  wire n3124;
  wire [33:0] n3125;
  wire [31:0] n3126;
  wire [31:0] n3128;
  wire [31:0] n3129;
  wire [33:0] n3130;
  wire n3131;
  wire n3133;
  wire n3134;
  wire [33:0] n3135;
  wire n3136;
  wire n3138;
  wire n3139;
  wire [33:0] n3140;
  wire [31:0] n3141;
  wire [31:0] n3143;
  wire [31:0] n3144;
  wire [33:0] n3145;
  wire n3146;
  wire n3148;
  wire n3149;
  wire [33:0] n3150;
  wire n3151;
  wire n3153;
  wire n3154;
  wire [33:0] n3155;
  wire [31:0] n3156;
  wire [31:0] n3158;
  wire [31:0] n3159;
  wire [33:0] n3160;
  wire n3161;
  wire n3163;
  wire n3164;
  wire [33:0] n3165;
  wire n3166;
  wire n3168;
  wire n3169;
  wire [33:0] n3170;
  wire [31:0] n3171;
  wire [31:0] n3173;
  wire [31:0] n3174;
  wire [33:0] n3175;
  wire n3176;
  wire n3178;
  wire n3179;
  wire [33:0] n3180;
  wire n3181;
  wire n3183;
  wire n3184;
  wire [33:0] n3185;
  wire [2559:0] n3188;
  wire [1087:0] n3189;
  assign \main_rsp_o_main_rsp_o[data]  = n2423; //(module output)
  assign \main_rsp_o_main_rsp_o[ack]  = n2424; //(module output)
  assign \main_rsp_o_main_rsp_o[err]  = n2425; //(module output)
  assign \dev_00_req_o_dev_00_req_o[addr]  = n2427; //(module output)
  assign \dev_00_req_o_dev_00_req_o[data]  = n2428; //(module output)
  assign \dev_00_req_o_dev_00_req_o[ben]  = n2429; //(module output)
  assign \dev_00_req_o_dev_00_req_o[stb]  = n2430; //(module output)
  assign \dev_00_req_o_dev_00_req_o[rw]  = n2431; //(module output)
  assign \dev_00_req_o_dev_00_req_o[src]  = n2432; //(module output)
  assign \dev_00_req_o_dev_00_req_o[priv]  = n2433; //(module output)
  assign \dev_00_req_o_dev_00_req_o[amo]  = n2434; //(module output)
  assign \dev_00_req_o_dev_00_req_o[amoop]  = n2435; //(module output)
  assign \dev_00_req_o_dev_00_req_o[fence]  = n2436; //(module output)
  assign \dev_00_req_o_dev_00_req_o[sleep]  = n2437; //(module output)
  assign \dev_00_req_o_dev_00_req_o[debug]  = n2438; //(module output)
  assign \dev_01_req_o_dev_01_req_o[addr]  = n2441; //(module output)
  assign \dev_01_req_o_dev_01_req_o[data]  = n2442; //(module output)
  assign \dev_01_req_o_dev_01_req_o[ben]  = n2443; //(module output)
  assign \dev_01_req_o_dev_01_req_o[stb]  = n2444; //(module output)
  assign \dev_01_req_o_dev_01_req_o[rw]  = n2445; //(module output)
  assign \dev_01_req_o_dev_01_req_o[src]  = n2446; //(module output)
  assign \dev_01_req_o_dev_01_req_o[priv]  = n2447; //(module output)
  assign \dev_01_req_o_dev_01_req_o[amo]  = n2448; //(module output)
  assign \dev_01_req_o_dev_01_req_o[amoop]  = n2449; //(module output)
  assign \dev_01_req_o_dev_01_req_o[fence]  = n2450; //(module output)
  assign \dev_01_req_o_dev_01_req_o[sleep]  = n2451; //(module output)
  assign \dev_01_req_o_dev_01_req_o[debug]  = n2452; //(module output)
  assign \dev_02_req_o_dev_02_req_o[addr]  = n2455; //(module output)
  assign \dev_02_req_o_dev_02_req_o[data]  = n2456; //(module output)
  assign \dev_02_req_o_dev_02_req_o[ben]  = n2457; //(module output)
  assign \dev_02_req_o_dev_02_req_o[stb]  = n2458; //(module output)
  assign \dev_02_req_o_dev_02_req_o[rw]  = n2459; //(module output)
  assign \dev_02_req_o_dev_02_req_o[src]  = n2460; //(module output)
  assign \dev_02_req_o_dev_02_req_o[priv]  = n2461; //(module output)
  assign \dev_02_req_o_dev_02_req_o[amo]  = n2462; //(module output)
  assign \dev_02_req_o_dev_02_req_o[amoop]  = n2463; //(module output)
  assign \dev_02_req_o_dev_02_req_o[fence]  = n2464; //(module output)
  assign \dev_02_req_o_dev_02_req_o[sleep]  = n2465; //(module output)
  assign \dev_02_req_o_dev_02_req_o[debug]  = n2466; //(module output)
  assign \dev_03_req_o_dev_03_req_o[addr]  = n2469; //(module output)
  assign \dev_03_req_o_dev_03_req_o[data]  = n2470; //(module output)
  assign \dev_03_req_o_dev_03_req_o[ben]  = n2471; //(module output)
  assign \dev_03_req_o_dev_03_req_o[stb]  = n2472; //(module output)
  assign \dev_03_req_o_dev_03_req_o[rw]  = n2473; //(module output)
  assign \dev_03_req_o_dev_03_req_o[src]  = n2474; //(module output)
  assign \dev_03_req_o_dev_03_req_o[priv]  = n2475; //(module output)
  assign \dev_03_req_o_dev_03_req_o[amo]  = n2476; //(module output)
  assign \dev_03_req_o_dev_03_req_o[amoop]  = n2477; //(module output)
  assign \dev_03_req_o_dev_03_req_o[fence]  = n2478; //(module output)
  assign \dev_03_req_o_dev_03_req_o[sleep]  = n2479; //(module output)
  assign \dev_03_req_o_dev_03_req_o[debug]  = n2480; //(module output)
  assign \dev_04_req_o_dev_04_req_o[addr]  = n2483; //(module output)
  assign \dev_04_req_o_dev_04_req_o[data]  = n2484; //(module output)
  assign \dev_04_req_o_dev_04_req_o[ben]  = n2485; //(module output)
  assign \dev_04_req_o_dev_04_req_o[stb]  = n2486; //(module output)
  assign \dev_04_req_o_dev_04_req_o[rw]  = n2487; //(module output)
  assign \dev_04_req_o_dev_04_req_o[src]  = n2488; //(module output)
  assign \dev_04_req_o_dev_04_req_o[priv]  = n2489; //(module output)
  assign \dev_04_req_o_dev_04_req_o[amo]  = n2490; //(module output)
  assign \dev_04_req_o_dev_04_req_o[amoop]  = n2491; //(module output)
  assign \dev_04_req_o_dev_04_req_o[fence]  = n2492; //(module output)
  assign \dev_04_req_o_dev_04_req_o[sleep]  = n2493; //(module output)
  assign \dev_04_req_o_dev_04_req_o[debug]  = n2494; //(module output)
  assign \dev_05_req_o_dev_05_req_o[addr]  = n2497; //(module output)
  assign \dev_05_req_o_dev_05_req_o[data]  = n2498; //(module output)
  assign \dev_05_req_o_dev_05_req_o[ben]  = n2499; //(module output)
  assign \dev_05_req_o_dev_05_req_o[stb]  = n2500; //(module output)
  assign \dev_05_req_o_dev_05_req_o[rw]  = n2501; //(module output)
  assign \dev_05_req_o_dev_05_req_o[src]  = n2502; //(module output)
  assign \dev_05_req_o_dev_05_req_o[priv]  = n2503; //(module output)
  assign \dev_05_req_o_dev_05_req_o[amo]  = n2504; //(module output)
  assign \dev_05_req_o_dev_05_req_o[amoop]  = n2505; //(module output)
  assign \dev_05_req_o_dev_05_req_o[fence]  = n2506; //(module output)
  assign \dev_05_req_o_dev_05_req_o[sleep]  = n2507; //(module output)
  assign \dev_05_req_o_dev_05_req_o[debug]  = n2508; //(module output)
  assign \dev_06_req_o_dev_06_req_o[addr]  = n2511; //(module output)
  assign \dev_06_req_o_dev_06_req_o[data]  = n2512; //(module output)
  assign \dev_06_req_o_dev_06_req_o[ben]  = n2513; //(module output)
  assign \dev_06_req_o_dev_06_req_o[stb]  = n2514; //(module output)
  assign \dev_06_req_o_dev_06_req_o[rw]  = n2515; //(module output)
  assign \dev_06_req_o_dev_06_req_o[src]  = n2516; //(module output)
  assign \dev_06_req_o_dev_06_req_o[priv]  = n2517; //(module output)
  assign \dev_06_req_o_dev_06_req_o[amo]  = n2518; //(module output)
  assign \dev_06_req_o_dev_06_req_o[amoop]  = n2519; //(module output)
  assign \dev_06_req_o_dev_06_req_o[fence]  = n2520; //(module output)
  assign \dev_06_req_o_dev_06_req_o[sleep]  = n2521; //(module output)
  assign \dev_06_req_o_dev_06_req_o[debug]  = n2522; //(module output)
  assign \dev_07_req_o_dev_07_req_o[addr]  = n2525; //(module output)
  assign \dev_07_req_o_dev_07_req_o[data]  = n2526; //(module output)
  assign \dev_07_req_o_dev_07_req_o[ben]  = n2527; //(module output)
  assign \dev_07_req_o_dev_07_req_o[stb]  = n2528; //(module output)
  assign \dev_07_req_o_dev_07_req_o[rw]  = n2529; //(module output)
  assign \dev_07_req_o_dev_07_req_o[src]  = n2530; //(module output)
  assign \dev_07_req_o_dev_07_req_o[priv]  = n2531; //(module output)
  assign \dev_07_req_o_dev_07_req_o[amo]  = n2532; //(module output)
  assign \dev_07_req_o_dev_07_req_o[amoop]  = n2533; //(module output)
  assign \dev_07_req_o_dev_07_req_o[fence]  = n2534; //(module output)
  assign \dev_07_req_o_dev_07_req_o[sleep]  = n2535; //(module output)
  assign \dev_07_req_o_dev_07_req_o[debug]  = n2536; //(module output)
  assign \dev_08_req_o_dev_08_req_o[addr]  = n2539; //(module output)
  assign \dev_08_req_o_dev_08_req_o[data]  = n2540; //(module output)
  assign \dev_08_req_o_dev_08_req_o[ben]  = n2541; //(module output)
  assign \dev_08_req_o_dev_08_req_o[stb]  = n2542; //(module output)
  assign \dev_08_req_o_dev_08_req_o[rw]  = n2543; //(module output)
  assign \dev_08_req_o_dev_08_req_o[src]  = n2544; //(module output)
  assign \dev_08_req_o_dev_08_req_o[priv]  = n2545; //(module output)
  assign \dev_08_req_o_dev_08_req_o[amo]  = n2546; //(module output)
  assign \dev_08_req_o_dev_08_req_o[amoop]  = n2547; //(module output)
  assign \dev_08_req_o_dev_08_req_o[fence]  = n2548; //(module output)
  assign \dev_08_req_o_dev_08_req_o[sleep]  = n2549; //(module output)
  assign \dev_08_req_o_dev_08_req_o[debug]  = n2550; //(module output)
  assign \dev_09_req_o_dev_09_req_o[addr]  = n2553; //(module output)
  assign \dev_09_req_o_dev_09_req_o[data]  = n2554; //(module output)
  assign \dev_09_req_o_dev_09_req_o[ben]  = n2555; //(module output)
  assign \dev_09_req_o_dev_09_req_o[stb]  = n2556; //(module output)
  assign \dev_09_req_o_dev_09_req_o[rw]  = n2557; //(module output)
  assign \dev_09_req_o_dev_09_req_o[src]  = n2558; //(module output)
  assign \dev_09_req_o_dev_09_req_o[priv]  = n2559; //(module output)
  assign \dev_09_req_o_dev_09_req_o[amo]  = n2560; //(module output)
  assign \dev_09_req_o_dev_09_req_o[amoop]  = n2561; //(module output)
  assign \dev_09_req_o_dev_09_req_o[fence]  = n2562; //(module output)
  assign \dev_09_req_o_dev_09_req_o[sleep]  = n2563; //(module output)
  assign \dev_09_req_o_dev_09_req_o[debug]  = n2564; //(module output)
  assign \dev_10_req_o_dev_10_req_o[addr]  = n2567; //(module output)
  assign \dev_10_req_o_dev_10_req_o[data]  = n2568; //(module output)
  assign \dev_10_req_o_dev_10_req_o[ben]  = n2569; //(module output)
  assign \dev_10_req_o_dev_10_req_o[stb]  = n2570; //(module output)
  assign \dev_10_req_o_dev_10_req_o[rw]  = n2571; //(module output)
  assign \dev_10_req_o_dev_10_req_o[src]  = n2572; //(module output)
  assign \dev_10_req_o_dev_10_req_o[priv]  = n2573; //(module output)
  assign \dev_10_req_o_dev_10_req_o[amo]  = n2574; //(module output)
  assign \dev_10_req_o_dev_10_req_o[amoop]  = n2575; //(module output)
  assign \dev_10_req_o_dev_10_req_o[fence]  = n2576; //(module output)
  assign \dev_10_req_o_dev_10_req_o[sleep]  = n2577; //(module output)
  assign \dev_10_req_o_dev_10_req_o[debug]  = n2578; //(module output)
  assign \dev_11_req_o_dev_11_req_o[addr]  = n2581; //(module output)
  assign \dev_11_req_o_dev_11_req_o[data]  = n2582; //(module output)
  assign \dev_11_req_o_dev_11_req_o[ben]  = n2583; //(module output)
  assign \dev_11_req_o_dev_11_req_o[stb]  = n2584; //(module output)
  assign \dev_11_req_o_dev_11_req_o[rw]  = n2585; //(module output)
  assign \dev_11_req_o_dev_11_req_o[src]  = n2586; //(module output)
  assign \dev_11_req_o_dev_11_req_o[priv]  = n2587; //(module output)
  assign \dev_11_req_o_dev_11_req_o[amo]  = n2588; //(module output)
  assign \dev_11_req_o_dev_11_req_o[amoop]  = n2589; //(module output)
  assign \dev_11_req_o_dev_11_req_o[fence]  = n2590; //(module output)
  assign \dev_11_req_o_dev_11_req_o[sleep]  = n2591; //(module output)
  assign \dev_11_req_o_dev_11_req_o[debug]  = n2592; //(module output)
  assign \dev_12_req_o_dev_12_req_o[addr]  = n2595; //(module output)
  assign \dev_12_req_o_dev_12_req_o[data]  = n2596; //(module output)
  assign \dev_12_req_o_dev_12_req_o[ben]  = n2597; //(module output)
  assign \dev_12_req_o_dev_12_req_o[stb]  = n2598; //(module output)
  assign \dev_12_req_o_dev_12_req_o[rw]  = n2599; //(module output)
  assign \dev_12_req_o_dev_12_req_o[src]  = n2600; //(module output)
  assign \dev_12_req_o_dev_12_req_o[priv]  = n2601; //(module output)
  assign \dev_12_req_o_dev_12_req_o[amo]  = n2602; //(module output)
  assign \dev_12_req_o_dev_12_req_o[amoop]  = n2603; //(module output)
  assign \dev_12_req_o_dev_12_req_o[fence]  = n2604; //(module output)
  assign \dev_12_req_o_dev_12_req_o[sleep]  = n2605; //(module output)
  assign \dev_12_req_o_dev_12_req_o[debug]  = n2606; //(module output)
  assign \dev_13_req_o_dev_13_req_o[addr]  = n2609; //(module output)
  assign \dev_13_req_o_dev_13_req_o[data]  = n2610; //(module output)
  assign \dev_13_req_o_dev_13_req_o[ben]  = n2611; //(module output)
  assign \dev_13_req_o_dev_13_req_o[stb]  = n2612; //(module output)
  assign \dev_13_req_o_dev_13_req_o[rw]  = n2613; //(module output)
  assign \dev_13_req_o_dev_13_req_o[src]  = n2614; //(module output)
  assign \dev_13_req_o_dev_13_req_o[priv]  = n2615; //(module output)
  assign \dev_13_req_o_dev_13_req_o[amo]  = n2616; //(module output)
  assign \dev_13_req_o_dev_13_req_o[amoop]  = n2617; //(module output)
  assign \dev_13_req_o_dev_13_req_o[fence]  = n2618; //(module output)
  assign \dev_13_req_o_dev_13_req_o[sleep]  = n2619; //(module output)
  assign \dev_13_req_o_dev_13_req_o[debug]  = n2620; //(module output)
  assign \dev_14_req_o_dev_14_req_o[addr]  = n2623; //(module output)
  assign \dev_14_req_o_dev_14_req_o[data]  = n2624; //(module output)
  assign \dev_14_req_o_dev_14_req_o[ben]  = n2625; //(module output)
  assign \dev_14_req_o_dev_14_req_o[stb]  = n2626; //(module output)
  assign \dev_14_req_o_dev_14_req_o[rw]  = n2627; //(module output)
  assign \dev_14_req_o_dev_14_req_o[src]  = n2628; //(module output)
  assign \dev_14_req_o_dev_14_req_o[priv]  = n2629; //(module output)
  assign \dev_14_req_o_dev_14_req_o[amo]  = n2630; //(module output)
  assign \dev_14_req_o_dev_14_req_o[amoop]  = n2631; //(module output)
  assign \dev_14_req_o_dev_14_req_o[fence]  = n2632; //(module output)
  assign \dev_14_req_o_dev_14_req_o[sleep]  = n2633; //(module output)
  assign \dev_14_req_o_dev_14_req_o[debug]  = n2634; //(module output)
  assign \dev_15_req_o_dev_15_req_o[addr]  = n2637; //(module output)
  assign \dev_15_req_o_dev_15_req_o[data]  = n2638; //(module output)
  assign \dev_15_req_o_dev_15_req_o[ben]  = n2639; //(module output)
  assign \dev_15_req_o_dev_15_req_o[stb]  = n2640; //(module output)
  assign \dev_15_req_o_dev_15_req_o[rw]  = n2641; //(module output)
  assign \dev_15_req_o_dev_15_req_o[src]  = n2642; //(module output)
  assign \dev_15_req_o_dev_15_req_o[priv]  = n2643; //(module output)
  assign \dev_15_req_o_dev_15_req_o[amo]  = n2644; //(module output)
  assign \dev_15_req_o_dev_15_req_o[amoop]  = n2645; //(module output)
  assign \dev_15_req_o_dev_15_req_o[fence]  = n2646; //(module output)
  assign \dev_15_req_o_dev_15_req_o[sleep]  = n2647; //(module output)
  assign \dev_15_req_o_dev_15_req_o[debug]  = n2648; //(module output)
  assign \dev_16_req_o_dev_16_req_o[addr]  = n2651; //(module output)
  assign \dev_16_req_o_dev_16_req_o[data]  = n2652; //(module output)
  assign \dev_16_req_o_dev_16_req_o[ben]  = n2653; //(module output)
  assign \dev_16_req_o_dev_16_req_o[stb]  = n2654; //(module output)
  assign \dev_16_req_o_dev_16_req_o[rw]  = n2655; //(module output)
  assign \dev_16_req_o_dev_16_req_o[src]  = n2656; //(module output)
  assign \dev_16_req_o_dev_16_req_o[priv]  = n2657; //(module output)
  assign \dev_16_req_o_dev_16_req_o[amo]  = n2658; //(module output)
  assign \dev_16_req_o_dev_16_req_o[amoop]  = n2659; //(module output)
  assign \dev_16_req_o_dev_16_req_o[fence]  = n2660; //(module output)
  assign \dev_16_req_o_dev_16_req_o[sleep]  = n2661; //(module output)
  assign \dev_16_req_o_dev_16_req_o[debug]  = n2662; //(module output)
  assign \dev_17_req_o_dev_17_req_o[addr]  = n2665; //(module output)
  assign \dev_17_req_o_dev_17_req_o[data]  = n2666; //(module output)
  assign \dev_17_req_o_dev_17_req_o[ben]  = n2667; //(module output)
  assign \dev_17_req_o_dev_17_req_o[stb]  = n2668; //(module output)
  assign \dev_17_req_o_dev_17_req_o[rw]  = n2669; //(module output)
  assign \dev_17_req_o_dev_17_req_o[src]  = n2670; //(module output)
  assign \dev_17_req_o_dev_17_req_o[priv]  = n2671; //(module output)
  assign \dev_17_req_o_dev_17_req_o[amo]  = n2672; //(module output)
  assign \dev_17_req_o_dev_17_req_o[amoop]  = n2673; //(module output)
  assign \dev_17_req_o_dev_17_req_o[fence]  = n2674; //(module output)
  assign \dev_17_req_o_dev_17_req_o[sleep]  = n2675; //(module output)
  assign \dev_17_req_o_dev_17_req_o[debug]  = n2676; //(module output)
  assign \dev_18_req_o_dev_18_req_o[addr]  = n2679; //(module output)
  assign \dev_18_req_o_dev_18_req_o[data]  = n2680; //(module output)
  assign \dev_18_req_o_dev_18_req_o[ben]  = n2681; //(module output)
  assign \dev_18_req_o_dev_18_req_o[stb]  = n2682; //(module output)
  assign \dev_18_req_o_dev_18_req_o[rw]  = n2683; //(module output)
  assign \dev_18_req_o_dev_18_req_o[src]  = n2684; //(module output)
  assign \dev_18_req_o_dev_18_req_o[priv]  = n2685; //(module output)
  assign \dev_18_req_o_dev_18_req_o[amo]  = n2686; //(module output)
  assign \dev_18_req_o_dev_18_req_o[amoop]  = n2687; //(module output)
  assign \dev_18_req_o_dev_18_req_o[fence]  = n2688; //(module output)
  assign \dev_18_req_o_dev_18_req_o[sleep]  = n2689; //(module output)
  assign \dev_18_req_o_dev_18_req_o[debug]  = n2690; //(module output)
  assign \dev_19_req_o_dev_19_req_o[addr]  = n2693; //(module output)
  assign \dev_19_req_o_dev_19_req_o[data]  = n2694; //(module output)
  assign \dev_19_req_o_dev_19_req_o[ben]  = n2695; //(module output)
  assign \dev_19_req_o_dev_19_req_o[stb]  = n2696; //(module output)
  assign \dev_19_req_o_dev_19_req_o[rw]  = n2697; //(module output)
  assign \dev_19_req_o_dev_19_req_o[src]  = n2698; //(module output)
  assign \dev_19_req_o_dev_19_req_o[priv]  = n2699; //(module output)
  assign \dev_19_req_o_dev_19_req_o[amo]  = n2700; //(module output)
  assign \dev_19_req_o_dev_19_req_o[amoop]  = n2701; //(module output)
  assign \dev_19_req_o_dev_19_req_o[fence]  = n2702; //(module output)
  assign \dev_19_req_o_dev_19_req_o[sleep]  = n2703; //(module output)
  assign \dev_19_req_o_dev_19_req_o[debug]  = n2704; //(module output)
  assign \dev_20_req_o_dev_20_req_o[addr]  = n2707; //(module output)
  assign \dev_20_req_o_dev_20_req_o[data]  = n2708; //(module output)
  assign \dev_20_req_o_dev_20_req_o[ben]  = n2709; //(module output)
  assign \dev_20_req_o_dev_20_req_o[stb]  = n2710; //(module output)
  assign \dev_20_req_o_dev_20_req_o[rw]  = n2711; //(module output)
  assign \dev_20_req_o_dev_20_req_o[src]  = n2712; //(module output)
  assign \dev_20_req_o_dev_20_req_o[priv]  = n2713; //(module output)
  assign \dev_20_req_o_dev_20_req_o[amo]  = n2714; //(module output)
  assign \dev_20_req_o_dev_20_req_o[amoop]  = n2715; //(module output)
  assign \dev_20_req_o_dev_20_req_o[fence]  = n2716; //(module output)
  assign \dev_20_req_o_dev_20_req_o[sleep]  = n2717; //(module output)
  assign \dev_20_req_o_dev_20_req_o[debug]  = n2718; //(module output)
  assign \dev_21_req_o_dev_21_req_o[addr]  = n2721; //(module output)
  assign \dev_21_req_o_dev_21_req_o[data]  = n2722; //(module output)
  assign \dev_21_req_o_dev_21_req_o[ben]  = n2723; //(module output)
  assign \dev_21_req_o_dev_21_req_o[stb]  = n2724; //(module output)
  assign \dev_21_req_o_dev_21_req_o[rw]  = n2725; //(module output)
  assign \dev_21_req_o_dev_21_req_o[src]  = n2726; //(module output)
  assign \dev_21_req_o_dev_21_req_o[priv]  = n2727; //(module output)
  assign \dev_21_req_o_dev_21_req_o[amo]  = n2728; //(module output)
  assign \dev_21_req_o_dev_21_req_o[amoop]  = n2729; //(module output)
  assign \dev_21_req_o_dev_21_req_o[fence]  = n2730; //(module output)
  assign \dev_21_req_o_dev_21_req_o[sleep]  = n2731; //(module output)
  assign \dev_21_req_o_dev_21_req_o[debug]  = n2732; //(module output)
  assign \dev_22_req_o_dev_22_req_o[addr]  = n2735; //(module output)
  assign \dev_22_req_o_dev_22_req_o[data]  = n2736; //(module output)
  assign \dev_22_req_o_dev_22_req_o[ben]  = n2737; //(module output)
  assign \dev_22_req_o_dev_22_req_o[stb]  = n2738; //(module output)
  assign \dev_22_req_o_dev_22_req_o[rw]  = n2739; //(module output)
  assign \dev_22_req_o_dev_22_req_o[src]  = n2740; //(module output)
  assign \dev_22_req_o_dev_22_req_o[priv]  = n2741; //(module output)
  assign \dev_22_req_o_dev_22_req_o[amo]  = n2742; //(module output)
  assign \dev_22_req_o_dev_22_req_o[amoop]  = n2743; //(module output)
  assign \dev_22_req_o_dev_22_req_o[fence]  = n2744; //(module output)
  assign \dev_22_req_o_dev_22_req_o[sleep]  = n2745; //(module output)
  assign \dev_22_req_o_dev_22_req_o[debug]  = n2746; //(module output)
  assign \dev_23_req_o_dev_23_req_o[addr]  = n2749; //(module output)
  assign \dev_23_req_o_dev_23_req_o[data]  = n2750; //(module output)
  assign \dev_23_req_o_dev_23_req_o[ben]  = n2751; //(module output)
  assign \dev_23_req_o_dev_23_req_o[stb]  = n2752; //(module output)
  assign \dev_23_req_o_dev_23_req_o[rw]  = n2753; //(module output)
  assign \dev_23_req_o_dev_23_req_o[src]  = n2754; //(module output)
  assign \dev_23_req_o_dev_23_req_o[priv]  = n2755; //(module output)
  assign \dev_23_req_o_dev_23_req_o[amo]  = n2756; //(module output)
  assign \dev_23_req_o_dev_23_req_o[amoop]  = n2757; //(module output)
  assign \dev_23_req_o_dev_23_req_o[fence]  = n2758; //(module output)
  assign \dev_23_req_o_dev_23_req_o[sleep]  = n2759; //(module output)
  assign \dev_23_req_o_dev_23_req_o[debug]  = n2760; //(module output)
  assign \dev_24_req_o_dev_24_req_o[addr]  = n2763; //(module output)
  assign \dev_24_req_o_dev_24_req_o[data]  = n2764; //(module output)
  assign \dev_24_req_o_dev_24_req_o[ben]  = n2765; //(module output)
  assign \dev_24_req_o_dev_24_req_o[stb]  = n2766; //(module output)
  assign \dev_24_req_o_dev_24_req_o[rw]  = n2767; //(module output)
  assign \dev_24_req_o_dev_24_req_o[src]  = n2768; //(module output)
  assign \dev_24_req_o_dev_24_req_o[priv]  = n2769; //(module output)
  assign \dev_24_req_o_dev_24_req_o[amo]  = n2770; //(module output)
  assign \dev_24_req_o_dev_24_req_o[amoop]  = n2771; //(module output)
  assign \dev_24_req_o_dev_24_req_o[fence]  = n2772; //(module output)
  assign \dev_24_req_o_dev_24_req_o[sleep]  = n2773; //(module output)
  assign \dev_24_req_o_dev_24_req_o[debug]  = n2774; //(module output)
  assign \dev_25_req_o_dev_25_req_o[addr]  = n2777; //(module output)
  assign \dev_25_req_o_dev_25_req_o[data]  = n2778; //(module output)
  assign \dev_25_req_o_dev_25_req_o[ben]  = n2779; //(module output)
  assign \dev_25_req_o_dev_25_req_o[stb]  = n2780; //(module output)
  assign \dev_25_req_o_dev_25_req_o[rw]  = n2781; //(module output)
  assign \dev_25_req_o_dev_25_req_o[src]  = n2782; //(module output)
  assign \dev_25_req_o_dev_25_req_o[priv]  = n2783; //(module output)
  assign \dev_25_req_o_dev_25_req_o[amo]  = n2784; //(module output)
  assign \dev_25_req_o_dev_25_req_o[amoop]  = n2785; //(module output)
  assign \dev_25_req_o_dev_25_req_o[fence]  = n2786; //(module output)
  assign \dev_25_req_o_dev_25_req_o[sleep]  = n2787; //(module output)
  assign \dev_25_req_o_dev_25_req_o[debug]  = n2788; //(module output)
  assign \dev_26_req_o_dev_26_req_o[addr]  = n2791; //(module output)
  assign \dev_26_req_o_dev_26_req_o[data]  = n2792; //(module output)
  assign \dev_26_req_o_dev_26_req_o[ben]  = n2793; //(module output)
  assign \dev_26_req_o_dev_26_req_o[stb]  = n2794; //(module output)
  assign \dev_26_req_o_dev_26_req_o[rw]  = n2795; //(module output)
  assign \dev_26_req_o_dev_26_req_o[src]  = n2796; //(module output)
  assign \dev_26_req_o_dev_26_req_o[priv]  = n2797; //(module output)
  assign \dev_26_req_o_dev_26_req_o[amo]  = n2798; //(module output)
  assign \dev_26_req_o_dev_26_req_o[amoop]  = n2799; //(module output)
  assign \dev_26_req_o_dev_26_req_o[fence]  = n2800; //(module output)
  assign \dev_26_req_o_dev_26_req_o[sleep]  = n2801; //(module output)
  assign \dev_26_req_o_dev_26_req_o[debug]  = n2802; //(module output)
  assign \dev_27_req_o_dev_27_req_o[addr]  = n2805; //(module output)
  assign \dev_27_req_o_dev_27_req_o[data]  = n2806; //(module output)
  assign \dev_27_req_o_dev_27_req_o[ben]  = n2807; //(module output)
  assign \dev_27_req_o_dev_27_req_o[stb]  = n2808; //(module output)
  assign \dev_27_req_o_dev_27_req_o[rw]  = n2809; //(module output)
  assign \dev_27_req_o_dev_27_req_o[src]  = n2810; //(module output)
  assign \dev_27_req_o_dev_27_req_o[priv]  = n2811; //(module output)
  assign \dev_27_req_o_dev_27_req_o[amo]  = n2812; //(module output)
  assign \dev_27_req_o_dev_27_req_o[amoop]  = n2813; //(module output)
  assign \dev_27_req_o_dev_27_req_o[fence]  = n2814; //(module output)
  assign \dev_27_req_o_dev_27_req_o[sleep]  = n2815; //(module output)
  assign \dev_27_req_o_dev_27_req_o[debug]  = n2816; //(module output)
  assign \dev_28_req_o_dev_28_req_o[addr]  = n2819; //(module output)
  assign \dev_28_req_o_dev_28_req_o[data]  = n2820; //(module output)
  assign \dev_28_req_o_dev_28_req_o[ben]  = n2821; //(module output)
  assign \dev_28_req_o_dev_28_req_o[stb]  = n2822; //(module output)
  assign \dev_28_req_o_dev_28_req_o[rw]  = n2823; //(module output)
  assign \dev_28_req_o_dev_28_req_o[src]  = n2824; //(module output)
  assign \dev_28_req_o_dev_28_req_o[priv]  = n2825; //(module output)
  assign \dev_28_req_o_dev_28_req_o[amo]  = n2826; //(module output)
  assign \dev_28_req_o_dev_28_req_o[amoop]  = n2827; //(module output)
  assign \dev_28_req_o_dev_28_req_o[fence]  = n2828; //(module output)
  assign \dev_28_req_o_dev_28_req_o[sleep]  = n2829; //(module output)
  assign \dev_28_req_o_dev_28_req_o[debug]  = n2830; //(module output)
  assign \dev_29_req_o_dev_29_req_o[addr]  = n2833; //(module output)
  assign \dev_29_req_o_dev_29_req_o[data]  = n2834; //(module output)
  assign \dev_29_req_o_dev_29_req_o[ben]  = n2835; //(module output)
  assign \dev_29_req_o_dev_29_req_o[stb]  = n2836; //(module output)
  assign \dev_29_req_o_dev_29_req_o[rw]  = n2837; //(module output)
  assign \dev_29_req_o_dev_29_req_o[src]  = n2838; //(module output)
  assign \dev_29_req_o_dev_29_req_o[priv]  = n2839; //(module output)
  assign \dev_29_req_o_dev_29_req_o[amo]  = n2840; //(module output)
  assign \dev_29_req_o_dev_29_req_o[amoop]  = n2841; //(module output)
  assign \dev_29_req_o_dev_29_req_o[fence]  = n2842; //(module output)
  assign \dev_29_req_o_dev_29_req_o[sleep]  = n2843; //(module output)
  assign \dev_29_req_o_dev_29_req_o[debug]  = n2844; //(module output)
  assign \dev_30_req_o_dev_30_req_o[addr]  = n2847; //(module output)
  assign \dev_30_req_o_dev_30_req_o[data]  = n2848; //(module output)
  assign \dev_30_req_o_dev_30_req_o[ben]  = n2849; //(module output)
  assign \dev_30_req_o_dev_30_req_o[stb]  = n2850; //(module output)
  assign \dev_30_req_o_dev_30_req_o[rw]  = n2851; //(module output)
  assign \dev_30_req_o_dev_30_req_o[src]  = n2852; //(module output)
  assign \dev_30_req_o_dev_30_req_o[priv]  = n2853; //(module output)
  assign \dev_30_req_o_dev_30_req_o[amo]  = n2854; //(module output)
  assign \dev_30_req_o_dev_30_req_o[amoop]  = n2855; //(module output)
  assign \dev_30_req_o_dev_30_req_o[fence]  = n2856; //(module output)
  assign \dev_30_req_o_dev_30_req_o[sleep]  = n2857; //(module output)
  assign \dev_30_req_o_dev_30_req_o[debug]  = n2858; //(module output)
  assign \dev_31_req_o_dev_31_req_o[addr]  = n2861; //(module output)
  assign \dev_31_req_o_dev_31_req_o[data]  = n2862; //(module output)
  assign \dev_31_req_o_dev_31_req_o[ben]  = n2863; //(module output)
  assign \dev_31_req_o_dev_31_req_o[stb]  = n2864; //(module output)
  assign \dev_31_req_o_dev_31_req_o[rw]  = n2865; //(module output)
  assign \dev_31_req_o_dev_31_req_o[src]  = n2866; //(module output)
  assign \dev_31_req_o_dev_31_req_o[priv]  = n2867; //(module output)
  assign \dev_31_req_o_dev_31_req_o[amo]  = n2868; //(module output)
  assign \dev_31_req_o_dev_31_req_o[amoop]  = n2869; //(module output)
  assign \dev_31_req_o_dev_31_req_o[fence]  = n2870; //(module output)
  assign \dev_31_req_o_dev_31_req_o[sleep]  = n2871; //(module output)
  assign \dev_31_req_o_dev_31_req_o[debug]  = n2872; //(module output)
  assign n2421 = {\main_req_i_main_req_i[debug] , \main_req_i_main_req_i[sleep] , \main_req_i_main_req_i[fence] , \main_req_i_main_req_i[amoop] , \main_req_i_main_req_i[amo] , \main_req_i_main_req_i[priv] , \main_req_i_main_req_i[src] , \main_req_i_main_req_i[rw] , \main_req_i_main_req_i[stb] , \main_req_i_main_req_i[ben] , \main_req_i_main_req_i[data] , \main_req_i_main_req_i[addr] };
  assign n2423 = neorv32_bus_reg_inst_n2874[31:0]; // extract
  assign n2424 = neorv32_bus_reg_inst_n2874[32]; // extract
  assign n2425 = neorv32_bus_reg_inst_n2874[33]; // extract
  assign n2427 = n2897[31:0]; // extract
  assign n2428 = n2897[63:32]; // extract
  assign n2429 = n2897[67:64]; // extract
  assign n2430 = n2897[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:76:3  */
  assign n2431 = n2897[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:78:5  */
  assign n2432 = n2897[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:78:5  */
  assign n2433 = n2897[71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:78:5  */
  assign n2434 = n2897[72]; // extract
  assign n2435 = n2897[76:73]; // extract
  assign n2436 = n2897[77]; // extract
  assign n2437 = n2897[78]; // extract
  assign n2438 = n2897[79]; // extract
  assign n2439 = {\dev_00_rsp_i_dev_00_rsp_i[err] , \dev_00_rsp_i_dev_00_rsp_i[ack] , \dev_00_rsp_i_dev_00_rsp_i[data] };
  assign n2441 = n2898[31:0]; // extract
  assign n2442 = n2898[63:32]; // extract
  assign n2443 = n2898[67:64]; // extract
  assign n2444 = n2898[68]; // extract
  assign n2445 = n2898[69]; // extract
  assign n2446 = n2898[70]; // extract
  assign n2447 = n2898[71]; // extract
  assign n2448 = n2898[72]; // extract
  assign n2449 = n2898[76:73]; // extract
  assign n2450 = n2898[77]; // extract
  assign n2451 = n2898[78]; // extract
  assign n2452 = n2898[79]; // extract
  assign n2453 = {\dev_01_rsp_i_dev_01_rsp_i[err] , \dev_01_rsp_i_dev_01_rsp_i[ack] , \dev_01_rsp_i_dev_01_rsp_i[data] };
  assign n2455 = n2899[31:0]; // extract
  assign n2456 = n2899[63:32]; // extract
  assign n2457 = n2899[67:64]; // extract
  assign n2458 = n2899[68]; // extract
  assign n2459 = n2899[69]; // extract
  assign n2460 = n2899[70]; // extract
  assign n2461 = n2899[71]; // extract
  assign n2462 = n2899[72]; // extract
  assign n2463 = n2899[76:73]; // extract
  assign n2464 = n2899[77]; // extract
  assign n2465 = n2899[78]; // extract
  assign n2466 = n2899[79]; // extract
  assign n2467 = {\dev_02_rsp_i_dev_02_rsp_i[err] , \dev_02_rsp_i_dev_02_rsp_i[ack] , \dev_02_rsp_i_dev_02_rsp_i[data] };
  assign n2469 = n2900[31:0]; // extract
  assign n2470 = n2900[63:32]; // extract
  assign n2471 = n2900[67:64]; // extract
  assign n2472 = n2900[68]; // extract
  assign n2473 = n2900[69]; // extract
  assign n2474 = n2900[70]; // extract
  assign n2475 = n2900[71]; // extract
  assign n2476 = n2900[72]; // extract
  assign n2477 = n2900[76:73]; // extract
  assign n2478 = n2900[77]; // extract
  assign n2479 = n2900[78]; // extract
  assign n2480 = n2900[79]; // extract
  assign n2481 = {\dev_03_rsp_i_dev_03_rsp_i[err] , \dev_03_rsp_i_dev_03_rsp_i[ack] , \dev_03_rsp_i_dev_03_rsp_i[data] };
  assign n2483 = n2901[31:0]; // extract
  assign n2484 = n2901[63:32]; // extract
  assign n2485 = n2901[67:64]; // extract
  assign n2486 = n2901[68]; // extract
  assign n2487 = n2901[69]; // extract
  assign n2488 = n2901[70]; // extract
  assign n2489 = n2901[71]; // extract
  assign n2490 = n2901[72]; // extract
  assign n2491 = n2901[76:73]; // extract
  assign n2492 = n2901[77]; // extract
  assign n2493 = n2901[78]; // extract
  assign n2494 = n2901[79]; // extract
  assign n2495 = {\dev_04_rsp_i_dev_04_rsp_i[err] , \dev_04_rsp_i_dev_04_rsp_i[ack] , \dev_04_rsp_i_dev_04_rsp_i[data] };
  assign n2497 = n2902[31:0]; // extract
  assign n2498 = n2902[63:32]; // extract
  assign n2499 = n2902[67:64]; // extract
  assign n2500 = n2902[68]; // extract
  assign n2501 = n2902[69]; // extract
  assign n2502 = n2902[70]; // extract
  assign n2503 = n2902[71]; // extract
  assign n2504 = n2902[72]; // extract
  assign n2505 = n2902[76:73]; // extract
  assign n2506 = n2902[77]; // extract
  assign n2507 = n2902[78]; // extract
  assign n2508 = n2902[79]; // extract
  assign n2509 = {\dev_05_rsp_i_dev_05_rsp_i[err] , \dev_05_rsp_i_dev_05_rsp_i[ack] , \dev_05_rsp_i_dev_05_rsp_i[data] };
  assign n2511 = n2903[31:0]; // extract
  assign n2512 = n2903[63:32]; // extract
  assign n2513 = n2903[67:64]; // extract
  assign n2514 = n2903[68]; // extract
  assign n2515 = n2903[69]; // extract
  assign n2516 = n2903[70]; // extract
  assign n2517 = n2903[71]; // extract
  assign n2518 = n2903[72]; // extract
  assign n2519 = n2903[76:73]; // extract
  assign n2520 = n2903[77]; // extract
  assign n2521 = n2903[78]; // extract
  assign n2522 = n2903[79]; // extract
  assign n2523 = {\dev_06_rsp_i_dev_06_rsp_i[err] , \dev_06_rsp_i_dev_06_rsp_i[ack] , \dev_06_rsp_i_dev_06_rsp_i[data] };
  assign n2525 = n2904[31:0]; // extract
  assign n2526 = n2904[63:32]; // extract
  assign n2527 = n2904[67:64]; // extract
  assign n2528 = n2904[68]; // extract
  assign n2529 = n2904[69]; // extract
  assign n2530 = n2904[70]; // extract
  assign n2531 = n2904[71]; // extract
  assign n2532 = n2904[72]; // extract
  assign n2533 = n2904[76:73]; // extract
  assign n2534 = n2904[77]; // extract
  assign n2535 = n2904[78]; // extract
  assign n2536 = n2904[79]; // extract
  assign n2537 = {\dev_07_rsp_i_dev_07_rsp_i[err] , \dev_07_rsp_i_dev_07_rsp_i[ack] , \dev_07_rsp_i_dev_07_rsp_i[data] };
  assign n2539 = n2905[31:0]; // extract
  assign n2540 = n2905[63:32]; // extract
  assign n2541 = n2905[67:64]; // extract
  assign n2542 = n2905[68]; // extract
  assign n2543 = n2905[69]; // extract
  assign n2544 = n2905[70]; // extract
  assign n2545 = n2905[71]; // extract
  assign n2546 = n2905[72]; // extract
  assign n2547 = n2905[76:73]; // extract
  assign n2548 = n2905[77]; // extract
  assign n2549 = n2905[78]; // extract
  assign n2550 = n2905[79]; // extract
  assign n2551 = {\dev_08_rsp_i_dev_08_rsp_i[err] , \dev_08_rsp_i_dev_08_rsp_i[ack] , \dev_08_rsp_i_dev_08_rsp_i[data] };
  assign n2553 = n2906[31:0]; // extract
  assign n2554 = n2906[63:32]; // extract
  assign n2555 = n2906[67:64]; // extract
  assign n2556 = n2906[68]; // extract
  assign n2557 = n2906[69]; // extract
  assign n2558 = n2906[70]; // extract
  assign n2559 = n2906[71]; // extract
  assign n2560 = n2906[72]; // extract
  assign n2561 = n2906[76:73]; // extract
  assign n2562 = n2906[77]; // extract
  assign n2563 = n2906[78]; // extract
  assign n2564 = n2906[79]; // extract
  assign n2565 = {\dev_09_rsp_i_dev_09_rsp_i[err] , \dev_09_rsp_i_dev_09_rsp_i[ack] , \dev_09_rsp_i_dev_09_rsp_i[data] };
  assign n2567 = n2907[31:0]; // extract
  assign n2568 = n2907[63:32]; // extract
  assign n2569 = n2907[67:64]; // extract
  assign n2570 = n2907[68]; // extract
  assign n2571 = n2907[69]; // extract
  assign n2572 = n2907[70]; // extract
  assign n2573 = n2907[71]; // extract
  assign n2574 = n2907[72]; // extract
  assign n2575 = n2907[76:73]; // extract
  assign n2576 = n2907[77]; // extract
  assign n2577 = n2907[78]; // extract
  assign n2578 = n2907[79]; // extract
  assign n2579 = {\dev_10_rsp_i_dev_10_rsp_i[err] , \dev_10_rsp_i_dev_10_rsp_i[ack] , \dev_10_rsp_i_dev_10_rsp_i[data] };
  assign n2581 = n2908[31:0]; // extract
  assign n2582 = n2908[63:32]; // extract
  assign n2583 = n2908[67:64]; // extract
  assign n2584 = n2908[68]; // extract
  assign n2585 = n2908[69]; // extract
  assign n2586 = n2908[70]; // extract
  assign n2587 = n2908[71]; // extract
  assign n2588 = n2908[72]; // extract
  assign n2589 = n2908[76:73]; // extract
  assign n2590 = n2908[77]; // extract
  assign n2591 = n2908[78]; // extract
  assign n2592 = n2908[79]; // extract
  assign n2593 = {\dev_11_rsp_i_dev_11_rsp_i[err] , \dev_11_rsp_i_dev_11_rsp_i[ack] , \dev_11_rsp_i_dev_11_rsp_i[data] };
  assign n2595 = n2909[31:0]; // extract
  assign n2596 = n2909[63:32]; // extract
  assign n2597 = n2909[67:64]; // extract
  assign n2598 = n2909[68]; // extract
  assign n2599 = n2909[69]; // extract
  assign n2600 = n2909[70]; // extract
  assign n2601 = n2909[71]; // extract
  assign n2602 = n2909[72]; // extract
  assign n2603 = n2909[76:73]; // extract
  assign n2604 = n2909[77]; // extract
  assign n2605 = n2909[78]; // extract
  assign n2606 = n2909[79]; // extract
  assign n2607 = {\dev_12_rsp_i_dev_12_rsp_i[err] , \dev_12_rsp_i_dev_12_rsp_i[ack] , \dev_12_rsp_i_dev_12_rsp_i[data] };
  assign n2609 = n2910[31:0]; // extract
  assign n2610 = n2910[63:32]; // extract
  assign n2611 = n2910[67:64]; // extract
  assign n2612 = n2910[68]; // extract
  assign n2613 = n2910[69]; // extract
  assign n2614 = n2910[70]; // extract
  assign n2615 = n2910[71]; // extract
  assign n2616 = n2910[72]; // extract
  assign n2617 = n2910[76:73]; // extract
  assign n2618 = n2910[77]; // extract
  assign n2619 = n2910[78]; // extract
  assign n2620 = n2910[79]; // extract
  assign n2621 = {\dev_13_rsp_i_dev_13_rsp_i[err] , \dev_13_rsp_i_dev_13_rsp_i[ack] , \dev_13_rsp_i_dev_13_rsp_i[data] };
  assign n2623 = n2911[31:0]; // extract
  assign n2624 = n2911[63:32]; // extract
  assign n2625 = n2911[67:64]; // extract
  assign n2626 = n2911[68]; // extract
  assign n2627 = n2911[69]; // extract
  assign n2628 = n2911[70]; // extract
  assign n2629 = n2911[71]; // extract
  assign n2630 = n2911[72]; // extract
  assign n2631 = n2911[76:73]; // extract
  assign n2632 = n2911[77]; // extract
  assign n2633 = n2911[78]; // extract
  assign n2634 = n2911[79]; // extract
  assign n2635 = {\dev_14_rsp_i_dev_14_rsp_i[err] , \dev_14_rsp_i_dev_14_rsp_i[ack] , \dev_14_rsp_i_dev_14_rsp_i[data] };
  assign n2637 = n2912[31:0]; // extract
  assign n2638 = n2912[63:32]; // extract
  assign n2639 = n2912[67:64]; // extract
  assign n2640 = n2912[68]; // extract
  assign n2641 = n2912[69]; // extract
  assign n2642 = n2912[70]; // extract
  assign n2643 = n2912[71]; // extract
  assign n2644 = n2912[72]; // extract
  assign n2645 = n2912[76:73]; // extract
  assign n2646 = n2912[77]; // extract
  assign n2647 = n2912[78]; // extract
  assign n2648 = n2912[79]; // extract
  assign n2649 = {\dev_15_rsp_i_dev_15_rsp_i[err] , \dev_15_rsp_i_dev_15_rsp_i[ack] , \dev_15_rsp_i_dev_15_rsp_i[data] };
  assign n2651 = n2913[31:0]; // extract
  assign n2652 = n2913[63:32]; // extract
  assign n2653 = n2913[67:64]; // extract
  assign n2654 = n2913[68]; // extract
  assign n2655 = n2913[69]; // extract
  assign n2656 = n2913[70]; // extract
  assign n2657 = n2913[71]; // extract
  assign n2658 = n2913[72]; // extract
  assign n2659 = n2913[76:73]; // extract
  assign n2660 = n2913[77]; // extract
  assign n2661 = n2913[78]; // extract
  assign n2662 = n2913[79]; // extract
  assign n2663 = {\dev_16_rsp_i_dev_16_rsp_i[err] , \dev_16_rsp_i_dev_16_rsp_i[ack] , \dev_16_rsp_i_dev_16_rsp_i[data] };
  assign n2665 = n2914[31:0]; // extract
  assign n2666 = n2914[63:32]; // extract
  assign n2667 = n2914[67:64]; // extract
  assign n2668 = n2914[68]; // extract
  assign n2669 = n2914[69]; // extract
  assign n2670 = n2914[70]; // extract
  assign n2671 = n2914[71]; // extract
  assign n2672 = n2914[72]; // extract
  assign n2673 = n2914[76:73]; // extract
  assign n2674 = n2914[77]; // extract
  assign n2675 = n2914[78]; // extract
  assign n2676 = n2914[79]; // extract
  assign n2677 = {\dev_17_rsp_i_dev_17_rsp_i[err] , \dev_17_rsp_i_dev_17_rsp_i[ack] , \dev_17_rsp_i_dev_17_rsp_i[data] };
  assign n2679 = n2915[31:0]; // extract
  assign n2680 = n2915[63:32]; // extract
  assign n2681 = n2915[67:64]; // extract
  assign n2682 = n2915[68]; // extract
  assign n2683 = n2915[69]; // extract
  assign n2684 = n2915[70]; // extract
  assign n2685 = n2915[71]; // extract
  assign n2686 = n2915[72]; // extract
  assign n2687 = n2915[76:73]; // extract
  assign n2688 = n2915[77]; // extract
  assign n2689 = n2915[78]; // extract
  assign n2690 = n2915[79]; // extract
  assign n2691 = {\dev_18_rsp_i_dev_18_rsp_i[err] , \dev_18_rsp_i_dev_18_rsp_i[ack] , \dev_18_rsp_i_dev_18_rsp_i[data] };
  assign n2693 = n2916[31:0]; // extract
  assign n2694 = n2916[63:32]; // extract
  assign n2695 = n2916[67:64]; // extract
  assign n2696 = n2916[68]; // extract
  assign n2697 = n2916[69]; // extract
  assign n2698 = n2916[70]; // extract
  assign n2699 = n2916[71]; // extract
  assign n2700 = n2916[72]; // extract
  assign n2701 = n2916[76:73]; // extract
  assign n2702 = n2916[77]; // extract
  assign n2703 = n2916[78]; // extract
  assign n2704 = n2916[79]; // extract
  assign n2705 = {\dev_19_rsp_i_dev_19_rsp_i[err] , \dev_19_rsp_i_dev_19_rsp_i[ack] , \dev_19_rsp_i_dev_19_rsp_i[data] };
  assign n2707 = n2917[31:0]; // extract
  assign n2708 = n2917[63:32]; // extract
  assign n2709 = n2917[67:64]; // extract
  assign n2710 = n2917[68]; // extract
  assign n2711 = n2917[69]; // extract
  assign n2712 = n2917[70]; // extract
  assign n2713 = n2917[71]; // extract
  assign n2714 = n2917[72]; // extract
  assign n2715 = n2917[76:73]; // extract
  assign n2716 = n2917[77]; // extract
  assign n2717 = n2917[78]; // extract
  assign n2718 = n2917[79]; // extract
  assign n2719 = {\dev_20_rsp_i_dev_20_rsp_i[err] , \dev_20_rsp_i_dev_20_rsp_i[ack] , \dev_20_rsp_i_dev_20_rsp_i[data] };
  assign n2721 = n2918[31:0]; // extract
  assign n2722 = n2918[63:32]; // extract
  assign n2723 = n2918[67:64]; // extract
  assign n2724 = n2918[68]; // extract
  assign n2725 = n2918[69]; // extract
  assign n2726 = n2918[70]; // extract
  assign n2727 = n2918[71]; // extract
  assign n2728 = n2918[72]; // extract
  assign n2729 = n2918[76:73]; // extract
  assign n2730 = n2918[77]; // extract
  assign n2731 = n2918[78]; // extract
  assign n2732 = n2918[79]; // extract
  assign n2733 = {\dev_21_rsp_i_dev_21_rsp_i[err] , \dev_21_rsp_i_dev_21_rsp_i[ack] , \dev_21_rsp_i_dev_21_rsp_i[data] };
  assign n2735 = n2919[31:0]; // extract
  assign n2736 = n2919[63:32]; // extract
  assign n2737 = n2919[67:64]; // extract
  assign n2738 = n2919[68]; // extract
  assign n2739 = n2919[69]; // extract
  assign n2740 = n2919[70]; // extract
  assign n2741 = n2919[71]; // extract
  assign n2742 = n2919[72]; // extract
  assign n2743 = n2919[76:73]; // extract
  assign n2744 = n2919[77]; // extract
  assign n2745 = n2919[78]; // extract
  assign n2746 = n2919[79]; // extract
  assign n2747 = {\dev_22_rsp_i_dev_22_rsp_i[err] , \dev_22_rsp_i_dev_22_rsp_i[ack] , \dev_22_rsp_i_dev_22_rsp_i[data] };
  assign n2749 = n2920[31:0]; // extract
  assign n2750 = n2920[63:32]; // extract
  assign n2751 = n2920[67:64]; // extract
  assign n2752 = n2920[68]; // extract
  assign n2753 = n2920[69]; // extract
  assign n2754 = n2920[70]; // extract
  assign n2755 = n2920[71]; // extract
  assign n2756 = n2920[72]; // extract
  assign n2757 = n2920[76:73]; // extract
  assign n2758 = n2920[77]; // extract
  assign n2759 = n2920[78]; // extract
  assign n2760 = n2920[79]; // extract
  assign n2761 = {\dev_23_rsp_i_dev_23_rsp_i[err] , \dev_23_rsp_i_dev_23_rsp_i[ack] , \dev_23_rsp_i_dev_23_rsp_i[data] };
  assign n2763 = n2921[31:0]; // extract
  assign n2764 = n2921[63:32]; // extract
  assign n2765 = n2921[67:64]; // extract
  assign n2766 = n2921[68]; // extract
  assign n2767 = n2921[69]; // extract
  assign n2768 = n2921[70]; // extract
  assign n2769 = n2921[71]; // extract
  assign n2770 = n2921[72]; // extract
  assign n2771 = n2921[76:73]; // extract
  assign n2772 = n2921[77]; // extract
  assign n2773 = n2921[78]; // extract
  assign n2774 = n2921[79]; // extract
  assign n2775 = {\dev_24_rsp_i_dev_24_rsp_i[err] , \dev_24_rsp_i_dev_24_rsp_i[ack] , \dev_24_rsp_i_dev_24_rsp_i[data] };
  assign n2777 = n2922[31:0]; // extract
  assign n2778 = n2922[63:32]; // extract
  assign n2779 = n2922[67:64]; // extract
  assign n2780 = n2922[68]; // extract
  assign n2781 = n2922[69]; // extract
  assign n2782 = n2922[70]; // extract
  assign n2783 = n2922[71]; // extract
  assign n2784 = n2922[72]; // extract
  assign n2785 = n2922[76:73]; // extract
  assign n2786 = n2922[77]; // extract
  assign n2787 = n2922[78]; // extract
  assign n2788 = n2922[79]; // extract
  assign n2789 = {\dev_25_rsp_i_dev_25_rsp_i[err] , \dev_25_rsp_i_dev_25_rsp_i[ack] , \dev_25_rsp_i_dev_25_rsp_i[data] };
  assign n2791 = n2923[31:0]; // extract
  assign n2792 = n2923[63:32]; // extract
  assign n2793 = n2923[67:64]; // extract
  assign n2794 = n2923[68]; // extract
  assign n2795 = n2923[69]; // extract
  assign n2796 = n2923[70]; // extract
  assign n2797 = n2923[71]; // extract
  assign n2798 = n2923[72]; // extract
  assign n2799 = n2923[76:73]; // extract
  assign n2800 = n2923[77]; // extract
  assign n2801 = n2923[78]; // extract
  assign n2802 = n2923[79]; // extract
  assign n2803 = {\dev_26_rsp_i_dev_26_rsp_i[err] , \dev_26_rsp_i_dev_26_rsp_i[ack] , \dev_26_rsp_i_dev_26_rsp_i[data] };
  assign n2805 = n2924[31:0]; // extract
  assign n2806 = n2924[63:32]; // extract
  assign n2807 = n2924[67:64]; // extract
  assign n2808 = n2924[68]; // extract
  assign n2809 = n2924[69]; // extract
  assign n2810 = n2924[70]; // extract
  assign n2811 = n2924[71]; // extract
  assign n2812 = n2924[72]; // extract
  assign n2813 = n2924[76:73]; // extract
  assign n2814 = n2924[77]; // extract
  assign n2815 = n2924[78]; // extract
  assign n2816 = n2924[79]; // extract
  assign n2817 = {\dev_27_rsp_i_dev_27_rsp_i[err] , \dev_27_rsp_i_dev_27_rsp_i[ack] , \dev_27_rsp_i_dev_27_rsp_i[data] };
  assign n2819 = n2925[31:0]; // extract
  assign n2820 = n2925[63:32]; // extract
  assign n2821 = n2925[67:64]; // extract
  assign n2822 = n2925[68]; // extract
  assign n2823 = n2925[69]; // extract
  assign n2824 = n2925[70]; // extract
  assign n2825 = n2925[71]; // extract
  assign n2826 = n2925[72]; // extract
  assign n2827 = n2925[76:73]; // extract
  assign n2828 = n2925[77]; // extract
  assign n2829 = n2925[78]; // extract
  assign n2830 = n2925[79]; // extract
  assign n2831 = {\dev_28_rsp_i_dev_28_rsp_i[err] , \dev_28_rsp_i_dev_28_rsp_i[ack] , \dev_28_rsp_i_dev_28_rsp_i[data] };
  assign n2833 = n2926[31:0]; // extract
  assign n2834 = n2926[63:32]; // extract
  assign n2835 = n2926[67:64]; // extract
  assign n2836 = n2926[68]; // extract
  assign n2837 = n2926[69]; // extract
  assign n2838 = n2926[70]; // extract
  assign n2839 = n2926[71]; // extract
  assign n2840 = n2926[72]; // extract
  assign n2841 = n2926[76:73]; // extract
  assign n2842 = n2926[77]; // extract
  assign n2843 = n2926[78]; // extract
  assign n2844 = n2926[79]; // extract
  assign n2845 = {\dev_29_rsp_i_dev_29_rsp_i[err] , \dev_29_rsp_i_dev_29_rsp_i[ack] , \dev_29_rsp_i_dev_29_rsp_i[data] };
  assign n2847 = n2927[31:0]; // extract
  assign n2848 = n2927[63:32]; // extract
  assign n2849 = n2927[67:64]; // extract
  assign n2850 = n2927[68]; // extract
  assign n2851 = n2927[69]; // extract
  assign n2852 = n2927[70]; // extract
  assign n2853 = n2927[71]; // extract
  assign n2854 = n2927[72]; // extract
  assign n2855 = n2927[76:73]; // extract
  assign n2856 = n2927[77]; // extract
  assign n2857 = n2927[78]; // extract
  assign n2858 = n2927[79]; // extract
  assign n2859 = {\dev_30_rsp_i_dev_30_rsp_i[err] , \dev_30_rsp_i_dev_30_rsp_i[ack] , \dev_30_rsp_i_dev_30_rsp_i[data] };
  assign n2861 = n2928[31:0]; // extract
  assign n2862 = n2928[63:32]; // extract
  assign n2863 = n2928[67:64]; // extract
  assign n2864 = n2928[68]; // extract
  assign n2865 = n2928[69]; // extract
  assign n2866 = n2928[70]; // extract
  assign n2867 = n2928[71]; // extract
  assign n2868 = n2928[72]; // extract
  assign n2869 = n2928[76:73]; // extract
  assign n2870 = n2928[77]; // extract
  assign n2871 = n2928[78]; // extract
  assign n2872 = n2928[79]; // extract
  assign n2873 = {\dev_31_rsp_i_dev_31_rsp_i[err] , \dev_31_rsp_i_dev_31_rsp_i[ack] , \dev_31_rsp_i_dev_31_rsp_i[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:631:10  */
  assign dev_req = n3188; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:632:10  */
  assign dev_rsp = n3189; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:635:10  */
  assign main_req = neorv32_bus_reg_inst_n2875; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:636:10  */
  assign main_rsp = n3185; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:653:21  */
  assign neorv32_bus_reg_inst_n2874 = n2888; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:654:21  */
  assign neorv32_bus_reg_inst_n2875 = n2890; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:642:3  */
  neorv32_bus_reg_9159cb8bcee7fcb95582f140960cdae72788d326 neorv32_bus_reg_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .\host_req_i_host_req_i[addr] (n2876),
    .\host_req_i_host_req_i[data] (n2877),
    .\host_req_i_host_req_i[ben] (n2878),
    .\host_req_i_host_req_i[stb] (n2879),
    .\host_req_i_host_req_i[rw] (n2880),
    .\host_req_i_host_req_i[src] (n2881),
    .\host_req_i_host_req_i[priv] (n2882),
    .\host_req_i_host_req_i[amo] (n2883),
    .\host_req_i_host_req_i[amoop] (n2884),
    .\host_req_i_host_req_i[fence] (n2885),
    .\host_req_i_host_req_i[sleep] (n2886),
    .\host_req_i_host_req_i[debug] (n2887),
    .\device_rsp_i_device_rsp_i[data] (n2892),
    .\device_rsp_i_device_rsp_i[ack] (n2893),
    .\device_rsp_i_device_rsp_i[err] (n2894),
    .\host_rsp_o_host_rsp_o[data] (\neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[data] ),
    .\host_rsp_o_host_rsp_o[ack] (\neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[ack] ),
    .\host_rsp_o_host_rsp_o[err] (\neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[err] ),
    .\device_req_o_device_req_o[addr] (\neorv32_bus_reg_inst.device_req_o_device_req_o[addr] ),
    .\device_req_o_device_req_o[data] (\neorv32_bus_reg_inst.device_req_o_device_req_o[data] ),
    .\device_req_o_device_req_o[ben] (\neorv32_bus_reg_inst.device_req_o_device_req_o[ben] ),
    .\device_req_o_device_req_o[stb] (\neorv32_bus_reg_inst.device_req_o_device_req_o[stb] ),
    .\device_req_o_device_req_o[rw] (\neorv32_bus_reg_inst.device_req_o_device_req_o[rw] ),
    .\device_req_o_device_req_o[src] (\neorv32_bus_reg_inst.device_req_o_device_req_o[src] ),
    .\device_req_o_device_req_o[priv] (\neorv32_bus_reg_inst.device_req_o_device_req_o[priv] ),
    .\device_req_o_device_req_o[amo] (\neorv32_bus_reg_inst.device_req_o_device_req_o[amo] ),
    .\device_req_o_device_req_o[amoop] (\neorv32_bus_reg_inst.device_req_o_device_req_o[amoop] ),
    .\device_req_o_device_req_o[fence] (\neorv32_bus_reg_inst.device_req_o_device_req_o[fence] ),
    .\device_req_o_device_req_o[sleep] (\neorv32_bus_reg_inst.device_req_o_device_req_o[sleep] ),
    .\device_req_o_device_req_o[debug] (\neorv32_bus_reg_inst.device_req_o_device_req_o[debug] ));
  assign n2876 = n2421[31:0]; // extract
  assign n2877 = n2421[63:32]; // extract
  assign n2878 = n2421[67:64]; // extract
  assign n2879 = n2421[68]; // extract
  assign n2880 = n2421[69]; // extract
  assign n2881 = n2421[70]; // extract
  assign n2882 = n2421[71]; // extract
  assign n2883 = n2421[72]; // extract
  assign n2884 = n2421[76:73]; // extract
  assign n2885 = n2421[77]; // extract
  assign n2886 = n2421[78]; // extract
  assign n2887 = n2421[79]; // extract
  assign n2888 = {\neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[err] , \neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[ack] , \neorv32_bus_reg_inst.host_rsp_o_host_rsp_o[data] };
  assign n2890 = {\neorv32_bus_reg_inst.device_req_o_device_req_o[debug] , \neorv32_bus_reg_inst.device_req_o_device_req_o[sleep] , \neorv32_bus_reg_inst.device_req_o_device_req_o[fence] , \neorv32_bus_reg_inst.device_req_o_device_req_o[amoop] , \neorv32_bus_reg_inst.device_req_o_device_req_o[amo] , \neorv32_bus_reg_inst.device_req_o_device_req_o[priv] , \neorv32_bus_reg_inst.device_req_o_device_req_o[src] , \neorv32_bus_reg_inst.device_req_o_device_req_o[rw] , \neorv32_bus_reg_inst.device_req_o_device_req_o[stb] , \neorv32_bus_reg_inst.device_req_o_device_req_o[ben] , \neorv32_bus_reg_inst.device_req_o_device_req_o[data] , \neorv32_bus_reg_inst.device_req_o_device_req_o[addr] };
  assign n2892 = main_rsp[31:0]; // extract
  assign n2893 = main_rsp[32]; // extract
  assign n2894 = main_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:661:26  */
  assign n2897 = dev_req[2559:2480]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:662:26  */
  assign n2898 = dev_req[2479:2400]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:663:26  */
  assign n2899 = dev_req[2399:2320]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:664:26  */
  assign n2900 = dev_req[2319:2240]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:665:26  */
  assign n2901 = dev_req[2239:2160]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:666:26  */
  assign n2902 = dev_req[2159:2080]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:667:26  */
  assign n2903 = dev_req[2079:2000]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:668:26  */
  assign n2904 = dev_req[1999:1920]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:669:26  */
  assign n2905 = dev_req[1919:1840]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:670:26  */
  assign n2906 = dev_req[1839:1760]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:671:26  */
  assign n2907 = dev_req[1759:1680]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:672:26  */
  assign n2908 = dev_req[1679:1600]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:673:26  */
  assign n2909 = dev_req[1599:1520]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:674:26  */
  assign n2910 = dev_req[1519:1440]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:675:26  */
  assign n2911 = dev_req[1439:1360]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:676:26  */
  assign n2912 = dev_req[1359:1280]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:677:26  */
  assign n2913 = dev_req[1279:1200]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:678:26  */
  assign n2914 = dev_req[1199:1120]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:679:26  */
  assign n2915 = dev_req[1119:1040]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:680:26  */
  assign n2916 = dev_req[1039:960]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:681:26  */
  assign n2917 = dev_req[959:880]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:682:26  */
  assign n2918 = dev_req[879:800]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:683:26  */
  assign n2919 = dev_req[799:720]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:684:26  */
  assign n2920 = dev_req[719:640]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:685:26  */
  assign n2921 = dev_req[639:560]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:686:26  */
  assign n2922 = dev_req[559:480]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:687:26  */
  assign n2923 = dev_req[479:400]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:688:26  */
  assign n2924 = dev_req[399:320]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:689:26  */
  assign n2925 = dev_req[319:240]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:690:26  */
  assign n2926 = dev_req[239:160]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:691:26  */
  assign n2927 = dev_req[159:80]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:692:26  */
  assign n2928 = dev_req[79:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n2930 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n2932 = n2930 == 5'b00000;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n2933 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n2935 = n2932 ? n2933 : 1'b0;
  assign n2936 = main_req[79:69]; // extract
  assign n2937 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n2941 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n2943 = n2941 == 5'b01111;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n2944 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n2946 = n2943 ? n2944 : 1'b0;
  assign n2947 = main_req[79:69]; // extract
  assign n2948 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n2951 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n2953 = n2951 == 5'b10000;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n2954 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n2956 = n2953 ? n2954 : 1'b0;
  assign n2957 = main_req[79:69]; // extract
  assign n2958 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n2961 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n2963 = n2961 == 5'b10100;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n2964 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n2966 = n2963 ? n2964 : 1'b0;
  assign n2967 = main_req[79:69]; // extract
  assign n2968 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n2971 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n2973 = n2971 == 5'b10101;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n2974 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n2976 = n2973 ? n2974 : 1'b0;
  assign n2977 = main_req[79:69]; // extract
  assign n2978 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n2981 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n2983 = n2981 == 5'b11000;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n2984 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n2986 = n2983 ? n2984 : 1'b0;
  assign n2987 = main_req[79:69]; // extract
  assign n2988 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n2991 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n2993 = n2991 == 5'b11001;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n2994 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n2996 = n2993 ? n2994 : 1'b0;
  assign n2997 = main_req[79:69]; // extract
  assign n2998 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n3001 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n3003 = n3001 == 5'b11100;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n3004 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n3006 = n3003 ? n3004 : 1'b0;
  assign n3007 = main_req[79:69]; // extract
  assign n3008 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n3011 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n3013 = n3011 == 5'b11110;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n3014 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n3016 = n3013 ? n3014 : 1'b0;
  assign n3017 = main_req[79:69]; // extract
  assign n3018 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:26  */
  assign n3021 = main_req[20:16]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:55  */
  assign n3023 = n3021 == 5'b11111;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:706:38  */
  assign n3024 = main_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:705:9  */
  assign n3026 = n3023 ? n3024 : 1'b0;
  assign n3027 = main_req[79:69]; // extract
  assign n3028 = main_req[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3033 = n3032[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3035 = dev_rsp[1085:1054]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3036 = n3033 | n3035;
  assign n3038 = n3037[33:32]; // extract
  assign n3039 = {n3038, n3036};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3040 = n3039[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3042 = dev_rsp[1086]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3043 = n3040 | n3042;
  assign n3044 = n3037[33]; // extract
  assign n3045 = {n3044, n3043, n3036};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3046 = n3045[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3048 = dev_rsp[1087]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3049 = n3046 | n3048;
  assign n3050 = {n3049, n3043, n3036};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3051 = n3050[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3053 = dev_rsp[575:544]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3054 = n3051 | n3053;
  assign n3055 = {n3049, n3043, n3054};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3056 = n3055[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3058 = dev_rsp[576]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3059 = n3056 | n3058;
  assign n3060 = {n3049, n3059, n3054};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3061 = n3060[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3063 = dev_rsp[577]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3064 = n3061 | n3063;
  assign n3065 = {n3064, n3059, n3054};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3066 = n3065[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3068 = dev_rsp[541:510]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3069 = n3066 | n3068;
  assign n3070 = {n3064, n3059, n3069};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3071 = n3070[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3073 = dev_rsp[542]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3074 = n3071 | n3073;
  assign n3075 = {n3064, n3074, n3069};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3076 = n3075[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3078 = dev_rsp[543]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3079 = n3076 | n3078;
  assign n3080 = {n3079, n3074, n3069};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3081 = n3080[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3083 = dev_rsp[405:374]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3084 = n3081 | n3083;
  assign n3085 = {n3079, n3074, n3084};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3086 = n3085[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3088 = dev_rsp[406]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3089 = n3086 | n3088;
  assign n3090 = {n3079, n3089, n3084};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3091 = n3090[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3093 = dev_rsp[407]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3094 = n3091 | n3093;
  assign n3095 = {n3094, n3089, n3084};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3096 = n3095[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3098 = dev_rsp[371:340]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3099 = n3096 | n3098;
  assign n3100 = {n3094, n3089, n3099};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3101 = n3100[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3103 = dev_rsp[372]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3104 = n3101 | n3103;
  assign n3105 = {n3094, n3104, n3099};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3106 = n3105[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3108 = dev_rsp[373]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3109 = n3106 | n3108;
  assign n3110 = {n3109, n3104, n3099};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3111 = n3110[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3113 = dev_rsp[269:238]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3114 = n3111 | n3113;
  assign n3115 = {n3109, n3104, n3114};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3116 = n3115[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3118 = dev_rsp[270]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3119 = n3116 | n3118;
  assign n3120 = {n3109, n3119, n3114};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3121 = n3120[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3123 = dev_rsp[271]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3124 = n3121 | n3123;
  assign n3125 = {n3124, n3119, n3114};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3126 = n3125[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3128 = dev_rsp[235:204]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3129 = n3126 | n3128;
  assign n3130 = {n3124, n3119, n3129};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3131 = n3130[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3133 = dev_rsp[236]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3134 = n3131 | n3133;
  assign n3135 = {n3124, n3134, n3129};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3136 = n3135[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3138 = dev_rsp[237]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3139 = n3136 | n3138;
  assign n3140 = {n3139, n3134, n3129};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3141 = n3140[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3143 = dev_rsp[133:102]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3144 = n3141 | n3143;
  assign n3145 = {n3139, n3134, n3144};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3146 = n3145[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3148 = dev_rsp[134]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3149 = n3146 | n3148;
  assign n3150 = {n3139, n3149, n3144};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3151 = n3150[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3153 = dev_rsp[135]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3154 = n3151 | n3153;
  assign n3155 = {n3154, n3149, n3144};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3156 = n3155[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3158 = dev_rsp[65:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3159 = n3156 | n3158;
  assign n3160 = {n3154, n3149, n3159};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3161 = n3160[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3163 = dev_rsp[66]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3164 = n3161 | n3163;
  assign n3165 = {n3154, n3164, n3159};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3166 = n3165[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3168 = dev_rsp[67]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3169 = n3166 | n3168;
  assign n3170 = {n3169, n3164, n3159};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:29  */
  assign n3171 = n3170[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:48  */
  assign n3173 = dev_rsp[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:729:34  */
  assign n3174 = n3171 | n3173;
  assign n3175 = {n3169, n3164, n3174};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:29  */
  assign n3176 = n3175[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:48  */
  assign n3178 = dev_rsp[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:730:34  */
  assign n3179 = n3176 | n3178;
  assign n3180 = {n3169, n3179, n3174};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:29  */
  assign n3181 = n3180[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:48  */
  assign n3183 = dev_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:731:34  */
  assign n3184 = n3181 | n3183;
  assign n3185 = {n3184, n3179, n3174};
  assign n3188 = {n2936, n2935, n2937, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, n2947, n2946, n2948, n2957, n2956, n2958, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, n2967, n2966, n2968, n2977, n2976, n2978, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, n2987, n2986, n2988, n2997, n2996, n2998, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, n3007, n3006, n3008, 80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, n3017, n3016, n3018, n3027, n3026, n3028};
  assign n3189 = {n2439, n2453, n2467, n2481, n2495, n2509, n2523, n2537, n2551, n2565, n2579, n2593, n2607, n2621, n2635, n2649, n2663, n2677, n2691, n2705, n2719, n2733, n2747, n2761, n2775, n2789, n2803, n2817, n2831, n2845, n2859, n2873};
endmodule

module neorv32_xbus_255_5ba93c9db0cff93f52b521d7420e43f6eda2784f
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   input  [31:0] xbus_dat_i,
   input  xbus_ack_i,
   input  xbus_err_i,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output [31:0] xbus_adr_o,
   output [31:0] xbus_dat_o,
   output [2:0] xbus_tag_o,
   output xbus_we_o,
   output [3:0] xbus_sel_o,
   output xbus_stb_o,
   output xbus_cyc_o);
  wire [79:0] n2318;
  wire [31:0] n2320;
  wire n2321;
  wire n2322;
  wire [79:0] bus_req;
  wire [33:0] bus_rsp;
  wire [1:0] pending;
  wire timeout;
  wire [8:0] timecnt;
  wire [31:0] \reg_stage_inst.host_rsp_o_host_rsp_o[data] ;
  wire \reg_stage_inst.host_rsp_o_host_rsp_o[ack] ;
  wire \reg_stage_inst.host_rsp_o_host_rsp_o[err] ;
  wire [31:0] \reg_stage_inst.device_req_o_device_req_o[addr] ;
  wire [31:0] \reg_stage_inst.device_req_o_device_req_o[data] ;
  wire [3:0] \reg_stage_inst.device_req_o_device_req_o[ben] ;
  wire \reg_stage_inst.device_req_o_device_req_o[stb] ;
  wire \reg_stage_inst.device_req_o_device_req_o[rw] ;
  wire \reg_stage_inst.device_req_o_device_req_o[src] ;
  wire \reg_stage_inst.device_req_o_device_req_o[priv] ;
  wire \reg_stage_inst.device_req_o_device_req_o[amo] ;
  wire [3:0] \reg_stage_inst.device_req_o_device_req_o[amoop] ;
  wire \reg_stage_inst.device_req_o_device_req_o[fence] ;
  wire \reg_stage_inst.device_req_o_device_req_o[sleep] ;
  wire \reg_stage_inst.device_req_o_device_req_o[debug] ;
  wire [31:0] n2330;
  wire [31:0] n2331;
  wire [3:0] n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire [3:0] n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire [33:0] n2342;
  wire [79:0] n2344;
  wire [31:0] n2346;
  wire n2347;
  wire n2348;
  wire n2350;
  wire [8:0] n2353;
  wire n2354;
  wire n2355;
  wire [1:0] n2357;
  wire n2359;
  wire [8:0] n2361;
  wire n2362;
  wire [1:0] n2364;
  wire [1:0] n2366;
  wire n2368;
  wire n2369;
  wire n2370;
  wire [1:0] n2373;
  wire [1:0] n2374;
  wire [1:0] n2375;
  reg [1:0] n2376;
  reg [8:0] n2378;
  wire n2380;
  wire n2382;
  wire n2385;
  wire [31:0] n2396;
  wire [31:0] n2397;
  wire n2398;
  wire [3:0] n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire [1:0] n2406;
  wire n2407;
  wire [2:0] n2408;
  wire n2409;
  wire [31:0] n2410;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire [33:0] n2417;
  reg [1:0] n2418;
  reg n2419;
  reg [8:0] n2420;
  assign \bus_rsp_o_bus_rsp_o[data]  = n2320; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n2321; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n2322; //(module output)
  assign xbus_adr_o = n2396; //(module output)
  assign xbus_dat_o = n2397; //(module output)
  assign xbus_tag_o = n2408; //(module output)
  assign xbus_we_o = n2398; //(module output)
  assign xbus_sel_o = n2399; //(module output)
  assign xbus_stb_o = n2400; //(module output)
  assign xbus_cyc_o = n2403; //(module output)
  assign n2318 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n2320 = n2342[31:0]; // extract
  assign n2321 = n2342[32]; // extract
  assign n2322 = n2342[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:47:10  */
  assign bus_req = n2344; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:48:10  */
  assign bus_rsp = n2417; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:51:10  */
  assign pending = n2418; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:52:10  */
  assign timeout = n2419; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:53:10  */
  assign timecnt = n2420; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:59:3  */
  neorv32_bus_reg_1489f923c4dca729178b3e3233458550d8dddf29 reg_stage_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .\host_req_i_host_req_i[addr] (n2330),
    .\host_req_i_host_req_i[data] (n2331),
    .\host_req_i_host_req_i[ben] (n2332),
    .\host_req_i_host_req_i[stb] (n2333),
    .\host_req_i_host_req_i[rw] (n2334),
    .\host_req_i_host_req_i[src] (n2335),
    .\host_req_i_host_req_i[priv] (n2336),
    .\host_req_i_host_req_i[amo] (n2337),
    .\host_req_i_host_req_i[amoop] (n2338),
    .\host_req_i_host_req_i[fence] (n2339),
    .\host_req_i_host_req_i[sleep] (n2340),
    .\host_req_i_host_req_i[debug] (n2341),
    .\device_rsp_i_device_rsp_i[data] (n2346),
    .\device_rsp_i_device_rsp_i[ack] (n2347),
    .\device_rsp_i_device_rsp_i[err] (n2348),
    .\host_rsp_o_host_rsp_o[data] (\reg_stage_inst.host_rsp_o_host_rsp_o[data] ),
    .\host_rsp_o_host_rsp_o[ack] (\reg_stage_inst.host_rsp_o_host_rsp_o[ack] ),
    .\host_rsp_o_host_rsp_o[err] (\reg_stage_inst.host_rsp_o_host_rsp_o[err] ),
    .\device_req_o_device_req_o[addr] (\reg_stage_inst.device_req_o_device_req_o[addr] ),
    .\device_req_o_device_req_o[data] (\reg_stage_inst.device_req_o_device_req_o[data] ),
    .\device_req_o_device_req_o[ben] (\reg_stage_inst.device_req_o_device_req_o[ben] ),
    .\device_req_o_device_req_o[stb] (\reg_stage_inst.device_req_o_device_req_o[stb] ),
    .\device_req_o_device_req_o[rw] (\reg_stage_inst.device_req_o_device_req_o[rw] ),
    .\device_req_o_device_req_o[src] (\reg_stage_inst.device_req_o_device_req_o[src] ),
    .\device_req_o_device_req_o[priv] (\reg_stage_inst.device_req_o_device_req_o[priv] ),
    .\device_req_o_device_req_o[amo] (\reg_stage_inst.device_req_o_device_req_o[amo] ),
    .\device_req_o_device_req_o[amoop] (\reg_stage_inst.device_req_o_device_req_o[amoop] ),
    .\device_req_o_device_req_o[fence] (\reg_stage_inst.device_req_o_device_req_o[fence] ),
    .\device_req_o_device_req_o[sleep] (\reg_stage_inst.device_req_o_device_req_o[sleep] ),
    .\device_req_o_device_req_o[debug] (\reg_stage_inst.device_req_o_device_req_o[debug] ));
  assign n2330 = n2318[31:0]; // extract
  assign n2331 = n2318[63:32]; // extract
  assign n2332 = n2318[67:64]; // extract
  assign n2333 = n2318[68]; // extract
  assign n2334 = n2318[69]; // extract
  assign n2335 = n2318[70]; // extract
  assign n2336 = n2318[71]; // extract
  assign n2337 = n2318[72]; // extract
  assign n2338 = n2318[76:73]; // extract
  assign n2339 = n2318[77]; // extract
  assign n2340 = n2318[78]; // extract
  assign n2341 = n2318[79]; // extract
  assign n2342 = {\reg_stage_inst.host_rsp_o_host_rsp_o[err] , \reg_stage_inst.host_rsp_o_host_rsp_o[ack] , \reg_stage_inst.host_rsp_o_host_rsp_o[data] };
  assign n2344 = {\reg_stage_inst.device_req_o_device_req_o[debug] , \reg_stage_inst.device_req_o_device_req_o[sleep] , \reg_stage_inst.device_req_o_device_req_o[fence] , \reg_stage_inst.device_req_o_device_req_o[amoop] , \reg_stage_inst.device_req_o_device_req_o[amo] , \reg_stage_inst.device_req_o_device_req_o[priv] , \reg_stage_inst.device_req_o_device_req_o[src] , \reg_stage_inst.device_req_o_device_req_o[rw] , \reg_stage_inst.device_req_o_device_req_o[stb] , \reg_stage_inst.device_req_o_device_req_o[ben] , \reg_stage_inst.device_req_o_device_req_o[data] , \reg_stage_inst.device_req_o_device_req_o[addr] };
  assign n2346 = bus_rsp[31:0]; // extract
  assign n2347 = bus_rsp[32]; // extract
  assign n2348 = bus_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:78:16  */
  assign n2350 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:89:58  */
  assign n2353 = timecnt + 9'b000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:90:33  */
  assign n2354 = xbus_ack_i | xbus_err_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:90:55  */
  assign n2355 = n2354 | timeout;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:90:11  */
  assign n2357 = n2355 ? 2'b00 : pending;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:87:9  */
  assign n2359 = pending == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:96:58  */
  assign n2361 = timecnt + 9'b000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:97:33  */
  assign n2362 = xbus_err_i | timeout;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:99:11  */
  assign n2364 = xbus_ack_i ? 2'b10 : pending;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:97:11  */
  assign n2366 = n2362 ? 2'b00 : n2364;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:94:9  */
  assign n2368 = pending == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:106:23  */
  assign n2369 = bus_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:107:25  */
  assign n2370 = bus_req[72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:107:13  */
  assign n2373 = n2370 ? 2'b11 : 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:106:11  */
  assign n2374 = n2369 ? n2373 : pending;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:144:30  */
  assign n2375 = {n2368, n2359};
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:85:7  */
  always @*
    case (n2375)
      2'b10: n2376 = n2366;
      2'b01: n2376 = n2357;
      default: n2376 = n2374;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:85:7  */
  always @*
    case (n2375)
      2'b10: n2378 = n2361;
      2'b01: n2378 = n2353;
      default: n2378 = 9'b000000000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:117:52  */
  assign n2380 = timecnt == 9'b011111111;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:117:29  */
  assign n2382 = n2380 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:117:7  */
  assign n2385 = n2382 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:132:25  */
  assign n2396 = bus_req[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:133:25  */
  assign n2397 = bus_req[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:134:25  */
  assign n2398 = bus_req[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:135:25  */
  assign n2399 = bus_req[67:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:136:25  */
  assign n2400 = bus_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:137:25  */
  assign n2401 = bus_req[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:137:39  */
  assign n2402 = pending[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:137:29  */
  assign n2403 = n2401 | n2402;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:138:25  */
  assign n2404 = bus_req[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:138:29  */
  assign n2406 = {n2404, 1'b0};
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:138:45  */
  assign n2407 = bus_req[71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:138:35  */
  assign n2408 = {n2406, n2407};
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:141:43  */
  assign n2409 = pending[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:141:30  */
  assign n2410 = n2409 ? xbus_dat_i : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:142:26  */
  assign n2412 = pending[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:142:30  */
  assign n2413 = n2412 & xbus_ack_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:143:26  */
  assign n2414 = pending[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:143:46  */
  assign n2415 = xbus_err_i | timeout;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:143:30  */
  assign n2416 = n2414 & n2415;
  assign n2417 = {n2416, n2413, n2410};
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:82:5  */
  always @(posedge clk_i or posedge n2350)
    if (n2350)
      n2418 <= 2'b00;
    else
      n2418 <= n2376;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:82:5  */
  always @(posedge clk_i or posedge n2350)
    if (n2350)
      n2419 <= 1'b0;
    else
      n2419 <= n2385;
  /* ../../ext/neorv32/rtl/core/neorv32_xbus.vhd:82:5  */
  always @(posedge clk_i or posedge n2350)
    if (n2350)
      n2420 <= 9'b000000000;
    else
      n2420 <= n2378;
endmodule

module neorv32_cache_16_64_69f24bf1e9d58f38577f662be0ab41a8f51212bb
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \host_req_i_host_req_i[addr] ,
   input  [31:0] \host_req_i_host_req_i[data] ,
   input  [3:0] \host_req_i_host_req_i[ben] ,
   input  \host_req_i_host_req_i[stb] ,
   input  \host_req_i_host_req_i[rw] ,
   input  \host_req_i_host_req_i[src] ,
   input  \host_req_i_host_req_i[priv] ,
   input  \host_req_i_host_req_i[amo] ,
   input  [3:0] \host_req_i_host_req_i[amoop] ,
   input  \host_req_i_host_req_i[fence] ,
   input  \host_req_i_host_req_i[sleep] ,
   input  \host_req_i_host_req_i[debug] ,
   input  [31:0] \bus_rsp_i_bus_rsp_i[data] ,
   input  \bus_rsp_i_bus_rsp_i[ack] ,
   input  \bus_rsp_i_bus_rsp_i[err] ,
   output [31:0] \host_rsp_o_host_rsp_o[data] ,
   output \host_rsp_o_host_rsp_o[ack] ,
   output \host_rsp_o_host_rsp_o[err] ,
   output [31:0] \bus_req_o_bus_req_o[addr] ,
   output [31:0] \bus_req_o_bus_req_o[data] ,
   output [3:0] \bus_req_o_bus_req_o[ben] ,
   output \bus_req_o_bus_req_o[stb] ,
   output \bus_req_o_bus_req_o[rw] ,
   output \bus_req_o_bus_req_o[src] ,
   output \bus_req_o_bus_req_o[priv] ,
   output \bus_req_o_bus_req_o[amo] ,
   output [3:0] \bus_req_o_bus_req_o[amoop] ,
   output \bus_req_o_bus_req_o[fence] ,
   output \bus_req_o_bus_req_o[sleep] ,
   output \bus_req_o_bus_req_o[debug] );
  wire [79:0] n2164;
  wire [31:0] n2166;
  wire n2167;
  wire n2168;
  wire [31:0] n2170;
  wire [31:0] n2171;
  wire [3:0] n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire [3:0] n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire [33:0] n2182;
  wire dir_acc_d;
  wire [79:0] bus_req;
  wire [79:0] cache_req;
  wire [33:0] bus_rsp;
  wire [33:0] cache_rsp;
  wire [69:0] cache_in_host;
  wire [69:0] cache_in_bus;
  wire [69:0] cache_in;
  wire [32:0] cache_out;
  wire cache_stat_dirty;
  wire cache_stat_hit;
  wire [31:0] cache_stat_base;
  wire cache_cmd_inval;
  wire cache_cmd_new;
  wire cache_cmd_dirty;
  wire bus_cmd_sync;
  wire bus_cmd_miss;
  wire bus_cmd_busy;
  wire n2185;
  wire n2195;
  wire n2196;
  wire n2197;
  wire [10:0] n2198;
  wire [67:0] n2199;
  wire [33:0] neorv32_cache_host_inst_n2202;
  wire neorv32_cache_host_inst_n2203;
  wire neorv32_cache_host_inst_n2204;
  wire neorv32_cache_host_inst_n2205;
  wire [31:0] neorv32_cache_host_inst_n2206;
  wire [3:0] neorv32_cache_host_inst_n2207;
  wire neorv32_cache_host_inst_n2208;
  wire [31:0] neorv32_cache_host_inst_n2209;
  wire neorv32_cache_host_inst_n2210;
  wire [31:0] n2211;
  wire n2212;
  wire [31:0] \neorv32_cache_host_inst.rsp_o_rsp_o[data] ;
  wire \neorv32_cache_host_inst.rsp_o_rsp_o[ack] ;
  wire \neorv32_cache_host_inst.rsp_o_rsp_o[err] ;
  wire [31:0] n2213;
  wire [31:0] n2214;
  wire [3:0] n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire [3:0] n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire [33:0] n2225;
  wire neorv32_cache_memory_inst_n2244;
  wire neorv32_cache_memory_inst_n2245;
  wire [31:0] neorv32_cache_memory_inst_n2246;
  wire [31:0] n2247;
  wire [3:0] n2248;
  wire n2249;
  wire [31:0] n2250;
  wire n2251;
  wire [31:0] neorv32_cache_memory_inst_n2252;
  wire neorv32_cache_memory_inst_n2253;
  wire n2264;
  wire [69:0] n2265;
  wire [79:0] neorv32_cache_bus_inst_n2266;
  wire neorv32_cache_bus_inst_n2267;
  wire neorv32_cache_bus_inst_n2268;
  wire neorv32_cache_bus_inst_n2269;
  wire [31:0] neorv32_cache_bus_inst_n2270;
  wire [3:0] neorv32_cache_bus_inst_n2271;
  wire neorv32_cache_bus_inst_n2272;
  wire [31:0] neorv32_cache_bus_inst_n2273;
  wire neorv32_cache_bus_inst_n2274;
  wire [31:0] n2275;
  wire [31:0] \neorv32_cache_bus_inst.bus_req_o_bus_req_o[addr] ;
  wire [31:0] \neorv32_cache_bus_inst.bus_req_o_bus_req_o[data] ;
  wire [3:0] \neorv32_cache_bus_inst.bus_req_o_bus_req_o[ben] ;
  wire \neorv32_cache_bus_inst.bus_req_o_bus_req_o[stb] ;
  wire \neorv32_cache_bus_inst.bus_req_o_bus_req_o[rw] ;
  wire \neorv32_cache_bus_inst.bus_req_o_bus_req_o[src] ;
  wire \neorv32_cache_bus_inst.bus_req_o_bus_req_o[priv] ;
  wire \neorv32_cache_bus_inst.bus_req_o_bus_req_o[amo] ;
  wire [3:0] \neorv32_cache_bus_inst.bus_req_o_bus_req_o[amoop] ;
  wire \neorv32_cache_bus_inst.bus_req_o_bus_req_o[fence] ;
  wire \neorv32_cache_bus_inst.bus_req_o_bus_req_o[sleep] ;
  wire \neorv32_cache_bus_inst.bus_req_o_bus_req_o[debug] ;
  wire [31:0] n2276;
  wire [31:0] n2277;
  wire [3:0] n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire [3:0] n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire [79:0] n2288;
  wire [31:0] n2290;
  wire n2291;
  wire n2292;
  wire [79:0] n2312;
  wire [69:0] n2315;
  wire [69:0] n2316;
  wire [32:0] n2317;
  assign \host_rsp_o_host_rsp_o[data]  = n2166; //(module output)
  assign \host_rsp_o_host_rsp_o[ack]  = n2167; //(module output)
  assign \host_rsp_o_host_rsp_o[err]  = n2168; //(module output)
  assign \bus_req_o_bus_req_o[addr]  = n2170; //(module output)
  assign \bus_req_o_bus_req_o[data]  = n2171; //(module output)
  assign \bus_req_o_bus_req_o[ben]  = n2172; //(module output)
  assign \bus_req_o_bus_req_o[stb]  = n2173; //(module output)
  assign \bus_req_o_bus_req_o[rw]  = n2174; //(module output)
  assign \bus_req_o_bus_req_o[src]  = n2175; //(module output)
  assign \bus_req_o_bus_req_o[priv]  = n2176; //(module output)
  assign \bus_req_o_bus_req_o[amo]  = n2177; //(module output)
  assign \bus_req_o_bus_req_o[amoop]  = n2178; //(module output)
  assign \bus_req_o_bus_req_o[fence]  = n2179; //(module output)
  assign \bus_req_o_bus_req_o[sleep]  = n2180; //(module output)
  assign \bus_req_o_bus_req_o[debug]  = n2181; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:352:23  */
  assign n2164 = {\host_req_i_host_req_i[debug] , \host_req_i_host_req_i[sleep] , \host_req_i_host_req_i[fence] , \host_req_i_host_req_i[amoop] , \host_req_i_host_req_i[amo] , \host_req_i_host_req_i[priv] , \host_req_i_host_req_i[src] , \host_req_i_host_req_i[rw] , \host_req_i_host_req_i[stb] , \host_req_i_host_req_i[ben] , \host_req_i_host_req_i[data] , \host_req_i_host_req_i[addr] };
  assign n2166 = cache_rsp[31:0]; // extract
  assign n2167 = cache_rsp[32]; // extract
  assign n2168 = cache_rsp[33]; // extract
  assign n2170 = bus_req[31:0]; // extract
  assign n2171 = bus_req[63:32]; // extract
  assign n2172 = bus_req[67:64]; // extract
  assign n2173 = bus_req[68]; // extract
  assign n2174 = bus_req[69]; // extract
  assign n2175 = bus_req[70]; // extract
  assign n2176 = bus_req[71]; // extract
  assign n2177 = bus_req[72]; // extract
  assign n2178 = bus_req[76:73]; // extract
  assign n2179 = bus_req[77]; // extract
  assign n2180 = bus_req[78]; // extract
  assign n2181 = bus_req[79]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:352:23  */
  assign n2182 = {\bus_rsp_i_bus_rsp_i[err] , \bus_rsp_i_bus_rsp_i[ack] , \bus_rsp_i_bus_rsp_i[data] };
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:141:10  */
  assign dir_acc_d = n2185; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:144:10  */
  assign bus_req = neorv32_cache_bus_inst_n2266; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:144:41  */
  assign cache_req = n2312; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:145:10  */
  assign bus_rsp = n2182; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:145:41  */
  assign cache_rsp = neorv32_cache_host_inst_n2202; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:155:10  */
  assign cache_in_host = n2315; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:155:25  */
  assign cache_in_bus = n2316; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:155:39  */
  assign cache_in = n2265; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:161:10  */
  assign cache_out = n2317; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:164:10  */
  assign cache_stat_dirty = neorv32_cache_memory_inst_n2245; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:164:28  */
  assign cache_stat_hit = neorv32_cache_memory_inst_n2244; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:165:10  */
  assign cache_stat_base = neorv32_cache_memory_inst_n2246; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:168:10  */
  assign cache_cmd_inval = neorv32_cache_bus_inst_n2268; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:168:27  */
  assign cache_cmd_new = neorv32_cache_bus_inst_n2269; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:168:42  */
  assign cache_cmd_dirty = neorv32_cache_host_inst_n2205; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:168:59  */
  assign bus_cmd_sync = neorv32_cache_host_inst_n2203; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:168:73  */
  assign bus_cmd_miss = neorv32_cache_host_inst_n2204; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:168:87  */
  assign bus_cmd_busy = neorv32_cache_bus_inst_n2267; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:174:20  */
  assign n2185 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:188:33  */
  assign n2195 = n2164[68]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:188:42  */
  assign n2196 = ~dir_acc_d;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:188:37  */
  assign n2197 = n2195 & n2196;
  assign n2198 = n2164[79:69]; // extract
  assign n2199 = n2164[67:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:238:19  */
  assign neorv32_cache_host_inst_n2202 = n2225; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:252:29  */
  assign n2211 = cache_out[31:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:253:29  */
  assign n2212 = cache_out[32]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:228:3  */
  neorv32_cache_host_bf8b4530d8d246dd74ac53a13471bba17941dff7 neorv32_cache_host_inst (
    .rstn_i(rstn_i),
    .clk_i(clk_i),
    .\req_i_req_i[addr] (n2213),
    .\req_i_req_i[data] (n2214),
    .\req_i_req_i[ben] (n2215),
    .\req_i_req_i[stb] (n2216),
    .\req_i_req_i[rw] (n2217),
    .\req_i_req_i[src] (n2218),
    .\req_i_req_i[priv] (n2219),
    .\req_i_req_i[amo] (n2220),
    .\req_i_req_i[amoop] (n2221),
    .\req_i_req_i[fence] (n2222),
    .\req_i_req_i[sleep] (n2223),
    .\req_i_req_i[debug] (n2224),
    .bus_busy_i(bus_cmd_busy),
    .hit_i(cache_stat_hit),
    .rdata_i(n2211),
    .rstat_i(n2212),
    .\rsp_o_rsp_o[data] (\neorv32_cache_host_inst.rsp_o_rsp_o[data] ),
    .\rsp_o_rsp_o[ack] (\neorv32_cache_host_inst.rsp_o_rsp_o[ack] ),
    .\rsp_o_rsp_o[err] (\neorv32_cache_host_inst.rsp_o_rsp_o[err] ),
    .bus_sync_o(neorv32_cache_host_inst_n2203),
    .bus_miss_o(neorv32_cache_host_inst_n2204),
    .dirty_o(neorv32_cache_host_inst_n2205),
    .addr_o(neorv32_cache_host_inst_n2206),
    .we_o(neorv32_cache_host_inst_n2207),
    .swe_o(neorv32_cache_host_inst_n2208),
    .wdata_o(neorv32_cache_host_inst_n2209),
    .wstat_o(neorv32_cache_host_inst_n2210));
  assign n2213 = cache_req[31:0]; // extract
  assign n2214 = cache_req[63:32]; // extract
  assign n2215 = cache_req[67:64]; // extract
  assign n2216 = cache_req[68]; // extract
  assign n2217 = cache_req[69]; // extract
  assign n2218 = cache_req[70]; // extract
  assign n2219 = cache_req[71]; // extract
  assign n2220 = cache_req[72]; // extract
  assign n2221 = cache_req[76:73]; // extract
  assign n2222 = cache_req[77]; // extract
  assign n2223 = cache_req[78]; // extract
  assign n2224 = cache_req[79]; // extract
  assign n2225 = {\neorv32_cache_host_inst.rsp_o_rsp_o[err] , \neorv32_cache_host_inst.rsp_o_rsp_o[ack] , \neorv32_cache_host_inst.rsp_o_rsp_o[data] };
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:278:26  */
  assign n2247 = cache_in[31:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:279:26  */
  assign n2248 = cache_in[35:32]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:280:26  */
  assign n2249 = cache_in[36]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:281:26  */
  assign n2250 = cache_in[68:37]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:282:26  */
  assign n2251 = cache_in[69]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:259:3  */
  neorv32_cache_memory_16_64_bf8b4530d8d246dd74ac53a13471bba17941dff7 neorv32_cache_memory_inst (
    .rstn_i(rstn_i),
    .clk_i(clk_i),
    .inval_i(cache_cmd_inval),
    .new_i(cache_cmd_new),
    .dirty_i(cache_cmd_dirty),
    .addr_i(n2247),
    .we_i(n2248),
    .swe_i(n2249),
    .wdata_i(n2250),
    .wstat_i(n2251),
    .hit_o(neorv32_cache_memory_inst_n2244),
    .dirty_o(neorv32_cache_memory_inst_n2245),
    .base_o(neorv32_cache_memory_inst_n2246),
    .rdata_o(neorv32_cache_memory_inst_n2252),
    .rstat_o(neorv32_cache_memory_inst_n2253));
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:288:48  */
  assign n2264 = ~bus_cmd_busy;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:288:29  */
  assign n2265 = n2264 ? cache_in_host : cache_in_bus;
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:306:19  */
  assign neorv32_cache_bus_inst_n2266 = n2288; // (signal)
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:323:29  */
  assign n2275 = cache_out[31:0]; // extract
  /* ../../src/hdl/sg13g2//neorv32_cache.vhd:293:3  */
  neorv32_cache_bus_16_64_bf8b4530d8d246dd74ac53a13471bba17941dff7 neorv32_cache_bus_inst (
    .rstn_i(rstn_i),
    .clk_i(clk_i),
    .\host_req_i_host_req_i[addr] (n2276),
    .\host_req_i_host_req_i[data] (n2277),
    .\host_req_i_host_req_i[ben] (n2278),
    .\host_req_i_host_req_i[stb] (n2279),
    .\host_req_i_host_req_i[rw] (n2280),
    .\host_req_i_host_req_i[src] (n2281),
    .\host_req_i_host_req_i[priv] (n2282),
    .\host_req_i_host_req_i[amo] (n2283),
    .\host_req_i_host_req_i[amoop] (n2284),
    .\host_req_i_host_req_i[fence] (n2285),
    .\host_req_i_host_req_i[sleep] (n2286),
    .\host_req_i_host_req_i[debug] (n2287),
    .\bus_rsp_i_bus_rsp_i[data] (n2290),
    .\bus_rsp_i_bus_rsp_i[ack] (n2291),
    .\bus_rsp_i_bus_rsp_i[err] (n2292),
    .cmd_sync_i(bus_cmd_sync),
    .cmd_miss_i(bus_cmd_miss),
    .dirty_i(cache_stat_dirty),
    .base_i(cache_stat_base),
    .rdata_i(n2275),
    .\bus_req_o_bus_req_o[addr] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[addr] ),
    .\bus_req_o_bus_req_o[data] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[data] ),
    .\bus_req_o_bus_req_o[ben] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[ben] ),
    .\bus_req_o_bus_req_o[stb] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[stb] ),
    .\bus_req_o_bus_req_o[rw] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[rw] ),
    .\bus_req_o_bus_req_o[src] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[src] ),
    .\bus_req_o_bus_req_o[priv] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[priv] ),
    .\bus_req_o_bus_req_o[amo] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[amo] ),
    .\bus_req_o_bus_req_o[amoop] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[amoop] ),
    .\bus_req_o_bus_req_o[fence] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[fence] ),
    .\bus_req_o_bus_req_o[sleep] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[sleep] ),
    .\bus_req_o_bus_req_o[debug] (\neorv32_cache_bus_inst.bus_req_o_bus_req_o[debug] ),
    .cmd_busy_o(neorv32_cache_bus_inst_n2267),
    .inval_o(neorv32_cache_bus_inst_n2268),
    .new_o(neorv32_cache_bus_inst_n2269),
    .addr_o(neorv32_cache_bus_inst_n2270),
    .we_o(neorv32_cache_bus_inst_n2271),
    .swe_o(neorv32_cache_bus_inst_n2272),
    .wdata_o(neorv32_cache_bus_inst_n2273),
    .wstat_o(neorv32_cache_bus_inst_n2274));
  assign n2276 = n2164[31:0]; // extract
  assign n2277 = n2164[63:32]; // extract
  assign n2278 = n2164[67:64]; // extract
  assign n2279 = n2164[68]; // extract
  assign n2280 = n2164[69]; // extract
  assign n2281 = n2164[70]; // extract
  assign n2282 = n2164[71]; // extract
  assign n2283 = n2164[72]; // extract
  assign n2284 = n2164[76:73]; // extract
  assign n2285 = n2164[77]; // extract
  assign n2286 = n2164[78]; // extract
  assign n2287 = n2164[79]; // extract
  assign n2288 = {\neorv32_cache_bus_inst.bus_req_o_bus_req_o[debug] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[sleep] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[fence] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[amoop] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[amo] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[priv] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[src] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[rw] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[stb] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[ben] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[data] , \neorv32_cache_bus_inst.bus_req_o_bus_req_o[addr] };
  assign n2290 = bus_rsp[31:0]; // extract
  assign n2291 = bus_rsp[32]; // extract
  assign n2292 = bus_rsp[33]; // extract
  assign n2312 = {n2198, n2197, n2199};
  assign n2315 = {neorv32_cache_host_inst_n2210, neorv32_cache_host_inst_n2209, neorv32_cache_host_inst_n2208, neorv32_cache_host_inst_n2207, neorv32_cache_host_inst_n2206};
  assign n2316 = {neorv32_cache_bus_inst_n2274, neorv32_cache_bus_inst_n2273, neorv32_cache_bus_inst_n2272, neorv32_cache_bus_inst_n2271, neorv32_cache_bus_inst_n2270};
  assign n2317 = {neorv32_cache_memory_inst_n2253, neorv32_cache_memory_inst_n2252};
endmodule

module neorv32_xip_bf8b4530d8d246dd74ac53a13471bba17941dff7
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   input  [31:0] \xip_req_i_xip_req_i[addr] ,
   input  [31:0] \xip_req_i_xip_req_i[data] ,
   input  [3:0] \xip_req_i_xip_req_i[ben] ,
   input  \xip_req_i_xip_req_i[stb] ,
   input  \xip_req_i_xip_req_i[rw] ,
   input  \xip_req_i_xip_req_i[src] ,
   input  \xip_req_i_xip_req_i[priv] ,
   input  \xip_req_i_xip_req_i[amo] ,
   input  [3:0] \xip_req_i_xip_req_i[amoop] ,
   input  \xip_req_i_xip_req_i[fence] ,
   input  \xip_req_i_xip_req_i[sleep] ,
   input  \xip_req_i_xip_req_i[debug] ,
   input  [7:0] clkgen_i,
   input  spi_dat_i,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] ,
   output [31:0] \xip_rsp_o_xip_rsp_o[data] ,
   output \xip_rsp_o_xip_rsp_o[ack] ,
   output \xip_rsp_o_xip_rsp_o[err] ,
   output clkgen_en_o,
   output spi_csn_o,
   output spi_clk_o,
   output spi_dat_o);
  wire [79:0] n1750;
  wire [31:0] n1752;
  wire n1753;
  wire n1754;
  wire [79:0] n1755;
  wire [31:0] n1757;
  wire n1758;
  wire n1759;
  wire [26:0] ctrl;
  wire [31:0] spi_data_lo;
  wire [31:0] spi_data_hi;
  wire spi_trigger;
  wire [31:0] xip_addr;
  wire [74:0] arbiter;
  wire [3:0] cdiv_cnt;
  wire spi_clk_en;
  wire [106:0] phy_if;
  wire n1765;
  wire n1767;
  localparam [31:0] n1769 = 32'b00000000000000000000000000000000;
  wire n1770;
  wire n1771;
  wire [1:0] n1772;
  wire n1774;
  wire n1775;
  wire [2:0] n1776;
  wire n1777;
  wire n1778;
  wire [3:0] n1779;
  wire n1780;
  wire [1:0] n1781;
  wire [7:0] n1782;
  wire n1783;
  wire n1784;
  wire [3:0] n1785;
  wire [26:0] n1786;
  wire [1:0] n1788;
  wire n1790;
  wire [31:0] n1791;
  wire [1:0] n1793;
  wire n1795;
  wire [31:0] n1796;
  wire n1800;
  wire [1:0] n1801;
  wire n1802;
  wire [2:0] n1803;
  wire n1804;
  wire n1805;
  wire [3:0] n1806;
  wire n1807;
  wire [1:0] n1808;
  wire [7:0] n1809;
  wire n1810;
  wire n1811;
  wire [3:0] n1812;
  wire n1813;
  wire n1814;
  wire n1816;
  wire [31:0] n1817;
  wire n1819;
  localparam [31:0] n1820 = 32'b00000000000000000000000000000000;
  wire [1:0] n1821;
  wire n1822;
  wire n1823;
  reg n1824;
  wire [2:0] n1825;
  wire [2:0] n1826;
  reg [2:0] n1827;
  wire n1828;
  wire n1829;
  reg n1830;
  wire n1831;
  wire n1832;
  reg n1833;
  wire [3:0] n1834;
  wire [3:0] n1835;
  reg [3:0] n1836;
  wire n1837;
  wire n1838;
  reg n1839;
  wire [1:0] n1840;
  wire [1:0] n1841;
  reg [1:0] n1842;
  wire [7:0] n1843;
  wire [7:0] n1844;
  reg [7:0] n1845;
  wire n1846;
  wire n1847;
  reg n1848;
  wire n1849;
  wire n1850;
  reg n1851;
  wire [3:0] n1852;
  wire [3:0] n1853;
  reg [3:0] n1854;
  wire [2:0] n1855;
  wire [2:0] n1856;
  wire [2:0] n1857;
  reg [2:0] n1858;
  wire n1859;
  wire n1860;
  reg n1861;
  wire n1862;
  wire n1863;
  reg n1864;
  wire [31:0] n1865;
  wire [31:0] n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1871;
  wire [31:0] n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1877;
  wire [33:0] n1879;
  wire [25:0] n1899;
  wire [1:0] n1901;
  wire [31:0] n1902;
  wire [7:0] n1903;
  wire [31:0] n1905;
  wire n1907;
  wire [31:0] n1908;
  wire [15:0] n1909;
  wire [31:0] n1911;
  wire n1913;
  wire [31:0] n1914;
  wire [23:0] n1915;
  wire [31:0] n1917;
  wire n1919;
  wire [31:0] n1920;
  wire [2:0] n1921;
  reg [31:0] n1922;
  wire n1926;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire [2:0] n1939;
  wire [2:0] n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire [31:0] n1945;
  wire [31:0] n1946;
  wire [31:0] n1947;
  wire [31:0] n1948;
  wire [31:0] n1950;
  wire [2:0] n1951;
  wire n1953;
  wire n1954;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire [2:0] n1962;
  wire n1964;
  wire n1965;
  wire n1967;
  wire n1968;
  wire [2:0] n1969;
  wire [2:0] n1971;
  wire [2:0] n1972;
  wire [2:0] n1973;
  wire [2:0] n1974;
  wire [64:0] n1975;
  wire [64:0] n1982;
  wire [2:0] n1988;
  wire n1991;
  wire n1993;
  wire n1996;
  wire [7:0] n1997;
  wire [39:0] n1998;
  wire [71:0] n2000;
  wire [2:0] n2001;
  wire [63:0] n2002;
  wire [71:0] n2004;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire [2:0] n2014;
  wire [2:0] n2015;
  wire n2017;
  wire [25:0] n2018;
  wire [25:0] n2019;
  wire n2020;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire [2:0] n2030;
  wire n2031;
  wire n2032;
  wire n2034;
  wire n2038;
  wire [7:0] n2047;
  wire [7:0] n2050;
  wire [7:0] n2052;
  wire [7:0] n2054;
  wire [31:0] n2055;
  wire n2056;
  wire n2057;
  wire n2060;
  wire [2:0] n2061;
  wire n2063;
  wire n2067;
  wire [5:0] n2069;
  reg [31:0] n2070;
  reg n2071;
  reg n2072;
  reg [2:0] n2073;
  reg n2074;
  reg n2075;
  reg [71:0] n2076;
  wire [2:0] n2079;
  wire n2081;
  wire [2:0] n2082;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2089;
  wire n2091;
  wire n2092;
  wire [2:0] n2093;
  wire n2097;
  wire n2098;
  wire [3:0] n2099;
  wire n2100;
  wire [3:0] n2102;
  wire [3:0] n2104;
  wire n2107;
  wire [3:0] n2108;
  wire n2110;
  wire [3:0] n2112;
  wire n2114;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire neorv32_xip_phy_inst_n2130;
  wire [3:0] n2131;
  wire [71:0] n2132;
  wire [31:0] neorv32_xip_phy_inst_n2133;
  wire neorv32_xip_phy_inst_n2134;
  wire neorv32_xip_phy_inst_n2135;
  wire neorv32_xip_phy_inst_n2136;
  wire [26:0] n2147;
  reg [26:0] n2148;
  wire [31:0] n2149;
  reg [31:0] n2150;
  wire [31:0] n2151;
  reg [31:0] n2152;
  reg n2153;
  reg [2:0] n2154;
  reg [64:0] n2155;
  reg [2:0] n2156;
  wire [74:0] n2157;
  reg [3:0] n2158;
  reg n2159;
  wire [106:0] n2160;
  reg [33:0] n2161;
  wire [33:0] n2162;
  wire n2163;
  assign \bus_rsp_o_bus_rsp_o[data]  = n1752; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n1753; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n1754; //(module output)
  assign \xip_rsp_o_xip_rsp_o[data]  = n1757; //(module output)
  assign \xip_rsp_o_xip_rsp_o[ack]  = n1758; //(module output)
  assign \xip_rsp_o_xip_rsp_o[err]  = n1759; //(module output)
  assign clkgen_en_o = n2123; //(module output)
  assign spi_csn_o = neorv32_xip_phy_inst_n2134; //(module output)
  assign spi_clk_o = neorv32_xip_phy_inst_n2135; //(module output)
  assign spi_dat_o = neorv32_xip_phy_inst_n2136; //(module output)
  assign n1750 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:111:5  */
  assign n1752 = n2161[31:0]; // extract
  assign n1753 = n2161[32]; // extract
  assign n1754 = n2161[33]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:109:3  */
  assign n1755 = {\xip_req_i_xip_req_i[debug] , \xip_req_i_xip_req_i[sleep] , \xip_req_i_xip_req_i[fence] , \xip_req_i_xip_req_i[amoop] , \xip_req_i_xip_req_i[amo] , \xip_req_i_xip_req_i[priv] , \xip_req_i_xip_req_i[src] , \xip_req_i_xip_req_i[rw] , \xip_req_i_xip_req_i[stb] , \xip_req_i_xip_req_i[ben] , \xip_req_i_xip_req_i[data] , \xip_req_i_xip_req_i[addr] };
  assign n1757 = n2162[31:0]; // extract
  assign n1758 = n2162[32]; // extract
  assign n1759 = n2162[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:67:10  */
  assign ctrl = n2148; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:70:10  */
  assign spi_data_lo = n2150; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:71:10  */
  assign spi_data_hi = n2152; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:72:10  */
  assign spi_trigger = n2153; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:75:10  */
  assign xip_addr = n1922; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:88:10  */
  assign arbiter = n2157; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:91:10  */
  assign cdiv_cnt = n2158; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:92:10  */
  assign spi_clk_en = n2159; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:129:10  */
  assign phy_if = n2160; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:137:16  */
  assign n1765 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:145:35  */
  assign n1767 = n1750[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:152:21  */
  assign n1770 = n1750[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:155:23  */
  assign n1771 = n1750[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:157:29  */
  assign n1772 = n1750[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:157:42  */
  assign n1774 = n1772 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:158:81  */
  assign n1775 = n1750[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:159:81  */
  assign n1776 = n1750[35:33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:160:81  */
  assign n1777 = n1750[36]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:161:81  */
  assign n1778 = n1750[37]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:162:81  */
  assign n1779 = n1750[41:38]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:163:81  */
  assign n1780 = n1750[42]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:164:81  */
  assign n1781 = n1750[44:43]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:165:81  */
  assign n1782 = n1750[52:45]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:166:81  */
  assign n1783 = n1750[53]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:167:81  */
  assign n1784 = n1750[54]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:168:81  */
  assign n1785 = n1750[58:55]; // extract
  assign n1786 = {n1785, n1784, n1783, n1782, n1781, n1780, n1779, n1778, n1777, n1776, n1775};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:171:29  */
  assign n1788 = n1750[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:171:42  */
  assign n1790 = n1788 == 2'b10;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:172:38  */
  assign n1791 = n1750[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:175:29  */
  assign n1793 = n1750[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:175:42  */
  assign n1795 = n1793 == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:176:38  */
  assign n1796 = n1750[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:175:11  */
  assign n1800 = n1795 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:30  */
  assign n1801 = n1750[3:2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:184:83  */
  assign n1802 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:185:83  */
  assign n1803 = ctrl[3:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:186:83  */
  assign n1804 = ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:187:83  */
  assign n1805 = ctrl[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:188:83  */
  assign n1806 = ctrl[9:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:189:83  */
  assign n1807 = ctrl[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:190:83  */
  assign n1808 = ctrl[12:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:191:83  */
  assign n1809 = ctrl[20:13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:192:83  */
  assign n1810 = ctrl[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:193:83  */
  assign n1811 = ctrl[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:194:83  */
  assign n1812 = ctrl[26:23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:196:57  */
  assign n1813 = phy_if[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:197:58  */
  assign n1814 = arbiter[71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:183:13  */
  assign n1816 = n1801 == 2'b00;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:199:40  */
  assign n1817 = phy_if[106:75]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:198:13  */
  assign n1819 = n1801 == 2'b10;
  assign n1821 = {n1819, n1816};
  assign n1822 = n1817[0]; // extract
  assign n1823 = n1820[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1824 = n1822;
      2'b01: n1824 = n1802;
      default: n1824 = n1823;
    endcase
  assign n1825 = n1817[3:1]; // extract
  assign n1826 = n1820[3:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1827 = n1825;
      2'b01: n1827 = n1803;
      default: n1827 = n1826;
    endcase
  assign n1828 = n1817[4]; // extract
  assign n1829 = n1820[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1830 = n1828;
      2'b01: n1830 = n1804;
      default: n1830 = n1829;
    endcase
  assign n1831 = n1817[5]; // extract
  assign n1832 = n1820[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1833 = n1831;
      2'b01: n1833 = n1805;
      default: n1833 = n1832;
    endcase
  assign n1834 = n1817[9:6]; // extract
  assign n1835 = n1820[9:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1836 = n1834;
      2'b01: n1836 = n1806;
      default: n1836 = n1835;
    endcase
  assign n1837 = n1817[10]; // extract
  assign n1838 = n1820[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1839 = n1837;
      2'b01: n1839 = n1807;
      default: n1839 = n1838;
    endcase
  assign n1840 = n1817[12:11]; // extract
  assign n1841 = n1820[12:11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1842 = n1840;
      2'b01: n1842 = n1808;
      default: n1842 = n1841;
    endcase
  assign n1843 = n1817[20:13]; // extract
  assign n1844 = n1820[20:13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1845 = n1843;
      2'b01: n1845 = n1809;
      default: n1845 = n1844;
    endcase
  assign n1846 = n1817[21]; // extract
  assign n1847 = n1820[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1848 = n1846;
      2'b01: n1848 = n1810;
      default: n1848 = n1847;
    endcase
  assign n1849 = n1817[22]; // extract
  assign n1850 = n1820[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1851 = n1849;
      2'b01: n1851 = n1811;
      default: n1851 = n1850;
    endcase
  assign n1852 = n1817[26:23]; // extract
  assign n1853 = n1820[26:23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1854 = n1852;
      2'b01: n1854 = n1812;
      default: n1854 = n1853;
    endcase
  assign n1855 = n1817[29:27]; // extract
  assign n1856 = n1820[29:27]; // extract
  assign n1857 = n1769[29:27]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1858 = n1855;
      2'b01: n1858 = n1857;
      default: n1858 = n1856;
    endcase
  assign n1859 = n1817[30]; // extract
  assign n1860 = n1820[30]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1861 = n1859;
      2'b01: n1861 = n1813;
      default: n1861 = n1860;
    endcase
  assign n1862 = n1817[31]; // extract
  assign n1863 = n1820[31]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:182:11  */
  always @*
    case (n1821)
      2'b10: n1864 = n1862;
      2'b01: n1864 = n1814;
      default: n1864 = n1863;
    endcase
  assign n1865 = {n1864, n1861, n1858, n1854, n1851, n1848, n1845, n1842, n1839, n1836, n1833, n1830, n1827, n1824};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:155:9  */
  assign n1866 = n1771 ? 32'b00000000000000000000000000000000 : n1865;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:155:9  */
  assign n1867 = n1774 & n1771;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:155:9  */
  assign n1868 = n1790 & n1771;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:155:9  */
  assign n1869 = n1795 & n1771;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:155:9  */
  assign n1871 = n1771 ? n1800 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:152:7  */
  assign n1872 = n1770 ? n1866 : 32'b00000000000000000000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:152:7  */
  assign n1873 = n1867 & n1770;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:152:7  */
  assign n1874 = n1868 & n1770;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:152:7  */
  assign n1875 = n1869 & n1770;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:152:7  */
  assign n1877 = n1770 ? n1871 : 1'b0;
  assign n1879 = {1'b0, n1767, n1872};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:216:40  */
  assign n1899 = arbiter[33:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:218:14  */
  assign n1901 = ctrl[12:11]; // extract
  assign n1902 = {4'b0000, n1899, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:219:39  */
  assign n1903 = n1902[7:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:219:53  */
  assign n1905 = {n1903, 24'b000000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:219:7  */
  assign n1907 = n1901 == 2'b00;
  assign n1908 = {4'b0000, n1899, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:220:39  */
  assign n1909 = n1908[15:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:220:53  */
  assign n1911 = {n1909, 16'b0000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:220:7  */
  assign n1913 = n1901 == 2'b01;
  assign n1914 = {4'b0000, n1899, 2'b00};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:221:39  */
  assign n1915 = n1914[23:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:221:53  */
  assign n1917 = {n1915, 8'b00000000};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:221:7  */
  assign n1919 = n1901 == 2'b10;
  assign n1920 = {4'b0000, n1899, 2'b00};
  assign n1921 = {n1919, n1913, n1907};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:218:5  */
  always @*
    case (n1921)
      3'b100: n1922 = n1917;
      3'b010: n1922 = n1911;
      3'b001: n1922 = n1905;
      default: n1922 = n1920;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:231:16  */
  assign n1926 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:239:15  */
  assign n1933 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:239:31  */
  assign n1934 = ~n1933;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:239:46  */
  assign n1935 = ctrl[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:239:66  */
  assign n1936 = ~n1935;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:239:38  */
  assign n1937 = n1934 | n1936;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:242:34  */
  assign n1939 = arbiter[5:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:239:7  */
  assign n1940 = n1937 ? 3'b000 : n1939;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:245:21  */
  assign n1941 = n1755[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:245:47  */
  assign n1942 = n1755[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:245:50  */
  assign n1943 = ~n1942;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:245:32  */
  assign n1944 = n1943 & n1941;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:246:35  */
  assign n1945 = n1755[31:0]; // extract
  assign n1946 = arbiter[37:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:245:7  */
  assign n1947 = n1944 ? n1945 : n1946;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:248:68  */
  assign n1948 = arbiter[37:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:248:74  */
  assign n1950 = n1948 + 32'b00000000000000000000000000000100;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:250:19  */
  assign n1951 = arbiter[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:250:25  */
  assign n1953 = n1951 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:251:42  */
  assign n1954 = n1755[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:250:7  */
  assign n1956 = n1953 ? n1954 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:15  */
  assign n1957 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:31  */
  assign n1958 = ~n1957;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:46  */
  assign n1959 = ctrl[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:66  */
  assign n1960 = ~n1959;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:38  */
  assign n1961 = n1958 | n1960;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:85  */
  assign n1962 = arbiter[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:91  */
  assign n1964 = n1962 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:73  */
  assign n1965 = n1961 | n1964;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:258:29  */
  assign n1967 = arbiter[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:258:52  */
  assign n1968 = ~n1967;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:259:63  */
  assign n1969 = arbiter[74:72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:259:72  */
  assign n1971 = n1969 + 3'b001;
  assign n1972 = arbiter[74:72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:258:7  */
  assign n1973 = n1968 ? n1971 : n1972;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:256:7  */
  assign n1974 = n1965 ? 3'b000 : n1973;
  assign n1975 = {n1956, n1950, n1947};
  assign n1982 = {1'b0, 32'b00000000000000000000000000000000, 32'b00000000000000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:269:34  */
  assign n1988 = arbiter[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:274:31  */
  assign n1991 = arbiter[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:278:36  */
  assign n1993 = arbiter[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:278:59  */
  assign n1996 = n1993 | 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:279:25  */
  assign n1997 = ctrl[20:13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:279:64  */
  assign n1998 = {n1997, xip_addr};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:279:75  */
  assign n2000 = {n1998, 32'b00000000000000000000000000000000};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:282:18  */
  assign n2001 = arbiter[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:286:42  */
  assign n2002 = {spi_data_hi, spi_data_lo};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:286:56  */
  assign n2004 = {n2002, 8'b00000000};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:284:7  */
  assign n2008 = n2001 == 3'b000;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:293:23  */
  assign n2009 = n1755[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:294:25  */
  assign n2010 = n1755[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:294:28  */
  assign n2011 = ~n2010;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:294:11  */
  assign n2014 = n2011 ? 3'b010 : 3'b101;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:293:9  */
  assign n2015 = n2009 ? n2014 : n1988;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:291:7  */
  assign n2017 = n2001 == 3'b001;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:303:25  */
  assign n2018 = arbiter[33:8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:303:63  */
  assign n2019 = arbiter[65:40]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:303:39  */
  assign n2020 = n2018 == n2019;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:303:78  */
  assign n2022 = 1'b1 & n2020;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:304:28  */
  assign n2023 = arbiter[74]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:304:51  */
  assign n2024 = ~n2023;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:303:95  */
  assign n2025 = n2024 & n2022;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:303:9  */
  assign n2030 = n2025 ? 3'b100 : 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:303:9  */
  assign n2031 = n2025 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:303:9  */
  assign n2032 = n2025 ? n1996 : 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:301:7  */
  assign n2034 = n2001 == 3'b010;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:312:7  */
  assign n2038 = n2001 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1114:44  */
  assign n2047 = phy_if[106:99]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1114:44  */
  assign n2050 = phy_if[98:91]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1114:44  */
  assign n2052 = phy_if[90:83]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1114:44  */
  assign n2054 = phy_if[82:75]; // extract
  assign n2055 = {n2054, n2052, n2050, n2047};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:320:20  */
  assign n2056 = phy_if[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:320:25  */
  assign n2057 = ~n2056;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:320:9  */
  assign n2060 = n2057 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:320:9  */
  assign n2061 = n2057 ? 3'b001 : n1988;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:317:7  */
  assign n2063 = n2001 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:325:7  */
  assign n2067 = n2001 == 3'b101;
  assign n2069 = {n2067, n2063, n2038, n2034, n2017, n2008};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:282:5  */
  always @*
    case (n2069)
      6'b100000: n2070 = 32'b00000000000000000000000000000000;
      6'b010000: n2070 = n2055;
      6'b001000: n2070 = 32'b00000000000000000000000000000000;
      6'b000100: n2070 = 32'b00000000000000000000000000000000;
      6'b000010: n2070 = 32'b00000000000000000000000000000000;
      6'b000001: n2070 = 32'b00000000000000000000000000000000;
      default: n2070 = 32'b00000000000000000000000000000000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:282:5  */
  always @*
    case (n2069)
      6'b100000: n2071 = 1'b0;
      6'b010000: n2071 = n2060;
      6'b001000: n2071 = 1'b0;
      6'b000100: n2071 = 1'b0;
      6'b000010: n2071 = 1'b0;
      6'b000001: n2071 = 1'b0;
      default: n2071 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:282:5  */
  always @*
    case (n2069)
      6'b100000: n2072 = 1'b1;
      6'b010000: n2072 = n1991;
      6'b001000: n2072 = n1991;
      6'b000100: n2072 = n1991;
      6'b000010: n2072 = n1991;
      6'b000001: n2072 = n1991;
      default: n2072 = n1991;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:282:5  */
  always @*
    case (n2069)
      6'b100000: n2073 = 3'b001;
      6'b010000: n2073 = n2061;
      6'b001000: n2073 = 3'b100;
      6'b000100: n2073 = n2030;
      6'b000010: n2073 = n2015;
      6'b000001: n2073 = 3'b001;
      default: n2073 = 3'b001;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:282:5  */
  always @*
    case (n2069)
      6'b100000: n2074 = 1'b0;
      6'b010000: n2074 = 1'b0;
      6'b001000: n2074 = 1'b1;
      6'b000100: n2074 = n2031;
      6'b000010: n2074 = 1'b0;
      6'b000001: n2074 = spi_trigger;
      default: n2074 = 1'b0;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:282:5  */
  always @*
    case (n2069)
      6'b100000: n2075 = n1996;
      6'b010000: n2075 = n1996;
      6'b001000: n2075 = n1996;
      6'b000100: n2075 = n2032;
      6'b000010: n2075 = n1996;
      6'b000001: n2075 = 1'b1;
      default: n2075 = n1996;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:282:5  */
  always @*
    case (n2069)
      6'b100000: n2076 = n2000;
      6'b010000: n2076 = n2000;
      6'b001000: n2076 = n2000;
      6'b000100: n2076 = n2000;
      6'b000010: n2076 = n2000;
      6'b000001: n2076 = n2004;
      default: n2076 = n2000;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:338:37  */
  assign n2079 = arbiter[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:338:43  */
  assign n2081 = n2079 == 3'b011;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:338:65  */
  assign n2082 = arbiter[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:338:71  */
  assign n2084 = n2082 == 3'b100;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:338:53  */
  assign n2085 = n2081 | n2084;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:338:23  */
  assign n2086 = n2085 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:345:16  */
  assign n2089 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:350:15  */
  assign n2091 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:350:31  */
  assign n2092 = ~n2091;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:352:47  */
  assign n2093 = ctrl[3:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:353:18  */
  assign n2097 = ctrl[22]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:352:100  */
  assign n2098 = n2163 | n2097;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:354:28  */
  assign n2099 = ctrl[26:23]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:354:22  */
  assign n2100 = cdiv_cnt == n2099;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:358:60  */
  assign n2102 = cdiv_cnt + 4'b0001;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:354:9  */
  assign n2104 = n2100 ? 4'b0000 : n2102;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:354:9  */
  assign n2107 = n2100 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:352:7  */
  assign n2108 = n2098 ? n2104 : cdiv_cnt;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:352:7  */
  assign n2110 = n2098 ? n2107 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:350:7  */
  assign n2112 = n2092 ? 4'b0000 : n2108;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:350:7  */
  assign n2114 = n2092 ? 1'b0 : n2110;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:365:22  */
  assign n2123 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:377:25  */
  assign n2124 = ctrl[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:378:25  */
  assign n2125 = ctrl[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:379:25  */
  assign n2126 = ctrl[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:381:28  */
  assign n2127 = phy_if[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:382:28  */
  assign n2128 = phy_if[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:383:25  */
  assign n2129 = ctrl[21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:385:25  */
  assign n2131 = ctrl[9:6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:386:28  */
  assign n2132 = phy_if[74:3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:370:3  */
  neorv32_xip_phy neorv32_xip_phy_inst (
    .rstn_i(rstn_i),
    .clk_i(clk_i),
    .spi_clk_en_i(spi_clk_en),
    .cf_enable_i(n2124),
    .cf_cpha_i(n2125),
    .cf_cpol_i(n2126),
    .op_start_i(n2127),
    .op_final_i(n2128),
    .op_csen_i(n2129),
    .op_nbytes_i(n2131),
    .op_wdata_i(n2132),
    .spi_dat_i(spi_dat_i),
    .op_busy_o(neorv32_xip_phy_inst_n2130),
    .op_rdata_o(neorv32_xip_phy_inst_n2133),
    .spi_csn_o(neorv32_xip_phy_inst_n2134),
    .spi_clk_o(neorv32_xip_phy_inst_n2135),
    .spi_dat_o(neorv32_xip_phy_inst_n2136));
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:143:5  */
  assign n2147 = n1873 ? n1786 : ctrl;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:143:5  */
  always @(posedge clk_i or posedge n1765)
    if (n1765)
      n2148 <= 27'b000000000000000000000000000;
    else
      n2148 <= n2147;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:143:5  */
  assign n2149 = n1874 ? n1791 : spi_data_lo;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:143:5  */
  always @(posedge clk_i or posedge n1765)
    if (n1765)
      n2150 <= 32'b00000000000000000000000000000000;
    else
      n2150 <= n2149;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:143:5  */
  assign n2151 = n1875 ? n1796 : spi_data_hi;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:143:5  */
  always @(posedge clk_i or posedge n1765)
    if (n1765)
      n2152 <= 32'b00000000000000000000000000000000;
    else
      n2152 <= n2151;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:143:5  */
  always @(posedge clk_i or posedge n1765)
    if (n1765)
      n2153 <= 1'b0;
    else
      n2153 <= n1877;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:237:5  */
  always @(posedge clk_i or posedge n1926)
    if (n1926)
      n2154 <= 3'b000;
    else
      n2154 <= n1974;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:237:5  */
  always @(posedge clk_i or posedge n1926)
    if (n1926)
      n2155 <= n1982;
    else
      n2155 <= n1975;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:237:5  */
  always @(posedge clk_i or posedge n1926)
    if (n1926)
      n2156 <= 3'b000;
    else
      n2156 <= n1940;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:231:5  */
  assign n2157 = {n2154, n2086, n2155, n2073, n2156};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:348:5  */
  always @(posedge clk_i or posedge n2089)
    if (n2089)
      n2158 <= 4'b0000;
    else
      n2158 <= n2112;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:348:5  */
  always @(posedge clk_i or posedge n2089)
    if (n2089)
      n2159 <= 1'b0;
    else
      n2159 <= n2114;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:345:5  */
  assign n2160 = {neorv32_xip_phy_inst_n2133, n2076, neorv32_xip_phy_inst_n2130, n2075, n2074};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:143:5  */
  always @(posedge clk_i or posedge n1765)
    if (n1765)
      n2161 <= 34'b0000000000000000000000000000000000;
    else
      n2161 <= n1879;
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:137:5  */
  assign n2162 = {n2072, n2071, n2070};
  /* ../../ext/neorv32/rtl/core/neorv32_xip.vhd:352:23  */
  assign n2163 = clkgen_i[n2093 * 1 +: 1]; //(Bmux)
endmodule

module neorv32_dmem_16384
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \bus_req_i_bus_req_i[addr] ,
   input  [31:0] \bus_req_i_bus_req_i[data] ,
   input  [3:0] \bus_req_i_bus_req_i[ben] ,
   input  \bus_req_i_bus_req_i[stb] ,
   input  \bus_req_i_bus_req_i[rw] ,
   input  \bus_req_i_bus_req_i[src] ,
   input  \bus_req_i_bus_req_i[priv] ,
   input  \bus_req_i_bus_req_i[amo] ,
   input  [3:0] \bus_req_i_bus_req_i[amoop] ,
   input  \bus_req_i_bus_req_i[fence] ,
   input  \bus_req_i_bus_req_i[sleep] ,
   input  \bus_req_i_bus_req_i[debug] ,
   output [31:0] \bus_rsp_o_bus_rsp_o[data] ,
   output \bus_rsp_o_bus_rsp_o[ack] ,
   output \bus_rsp_o_bus_rsp_o[err] );
  wire [79:0] n1665;
  wire [31:0] n1667;
  wire n1668;
  wire n1669;
  wire [31:0] rdata;
  wire [31:0] wr_mask;
  wire rden;
  wire [11:0] addr;
  wire wen;
  wire ren;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire [15:0] \row_n1_inst.A_DOUT ;
  localparam n1677 = 1'b1;
  wire [15:0] n1678;
  localparam n1679 = 1'b1;
  wire [15:0] n1681;
  localparam n1682 = 1'b0;
  localparam n1683 = 1'b0;
  localparam n1684 = 1'b0;
  localparam n1685 = 1'b0;
  localparam n1686 = 1'b0;
  localparam [11:0] n1687 = 12'b000000000000;
  localparam [15:0] n1688 = 16'b0000000000000000;
  localparam [15:0] n1689 = 16'b0000000000000000;
  wire n1691;
  wire n1692;
  wire [7:0] n1693;
  wire n1696;
  wire n1697;
  wire [7:0] n1698;
  wire [15:0] \row_n2_inst.A_DOUT ;
  localparam n1700 = 1'b1;
  wire [15:0] n1701;
  localparam n1702 = 1'b1;
  wire [15:0] n1704;
  localparam n1705 = 1'b0;
  localparam n1706 = 1'b0;
  localparam n1707 = 1'b0;
  localparam n1708 = 1'b0;
  localparam n1709 = 1'b0;
  localparam [11:0] n1710 = 12'b000000000000;
  localparam [15:0] n1711 = 16'b0000000000000000;
  localparam [15:0] n1712 = 16'b0000000000000000;
  wire n1714;
  wire n1715;
  wire [7:0] n1716;
  wire n1719;
  wire n1720;
  wire [7:0] n1721;
  wire [11:0] n1724;
  wire n1726;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire [31:0] n1741;
  wire [31:0] n1744;
  wire [31:0] n1745;
  reg n1746;
  reg n1748;
  wire [33:0] n1749;
  assign \bus_rsp_o_bus_rsp_o[data]  = n1667; //(module output)
  assign \bus_rsp_o_bus_rsp_o[ack]  = n1668; //(module output)
  assign \bus_rsp_o_bus_rsp_o[err]  = n1669; //(module output)
  assign n1665 = {\bus_req_i_bus_req_i[debug] , \bus_req_i_bus_req_i[sleep] , \bus_req_i_bus_req_i[fence] , \bus_req_i_bus_req_i[amoop] , \bus_req_i_bus_req_i[amo] , \bus_req_i_bus_req_i[priv] , \bus_req_i_bus_req_i[src] , \bus_req_i_bus_req_i[rw] , \bus_req_i_bus_req_i[stb] , \bus_req_i_bus_req_i[ben] , \bus_req_i_bus_req_i[data] , \bus_req_i_bus_req_i[addr] };
  assign n1667 = n1749[31:0]; // extract
  assign n1668 = n1749[32]; // extract
  assign n1669 = n1749[33]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:39:10  */
  assign rdata = n1744; // (signal)
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:40:10  */
  assign wr_mask = n1745; // (signal)
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:41:10  */
  assign rden = n1746; // (signal)
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:42:10  */
  assign addr = n1724; // (signal)
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:44:10  */
  assign wen = n1672; // (signal)
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:44:15  */
  assign ren = n1676; // (signal)
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:74:20  */
  assign n1670 = n1665[68]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:74:38  */
  assign n1671 = n1665[69]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:74:24  */
  assign n1672 = n1670 & n1671;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:75:20  */
  assign n1673 = n1665[68]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:75:42  */
  assign n1674 = n1665[69]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:75:28  */
  assign n1675 = ~n1674;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:75:24  */
  assign n1676 = n1673 & n1675;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:79:5  */
  RM_IHPSG13_1P_4096x16_c3_bm_bist row_n1_inst (
    .A_CLK(clk_i),
    .A_MEN(n1677),
    .A_WEN(wen),
    .A_REN(ren),
    .A_ADDR(addr),
    .A_DIN(n1678),
    .A_DLY(n1679),
    .A_BM(n1681),
    .A_BIST_CLK(n1682),
    .A_BIST_EN(n1683),
    .A_BIST_MEN(n1684),
    .A_BIST_WEN(n1685),
    .A_BIST_REN(n1686),
    .A_BIST_ADDR(n1687),
    .A_BIST_DIN(n1688),
    .A_BIST_BM(n1689),
    .A_DOUT(\row_n1_inst.A_DOUT ));
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:86:49  */
  assign n1678 = n1665[47:32]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:89:24  */
  assign n1681 = wr_mask[15:0]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:99:60  */
  assign n1691 = n1665[64]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:99:66  */
  assign n1692 = ~n1691;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:99:42  */
  assign n1693 = n1692 ? 8'b00000000 : 8'b11111111;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:100:63  */
  assign n1696 = n1665[65]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:100:71  */
  assign n1697 = ~n1696;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:100:45  */
  assign n1698 = n1697 ? 8'b00000000 : 8'b11111111;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:79:5  */
  RM_IHPSG13_1P_4096x16_c3_bm_bist row_n2_inst (
    .A_CLK(clk_i),
    .A_MEN(n1700),
    .A_WEN(wen),
    .A_REN(ren),
    .A_ADDR(addr),
    .A_DIN(n1701),
    .A_DLY(n1702),
    .A_BM(n1704),
    .A_BIST_CLK(n1705),
    .A_BIST_EN(n1706),
    .A_BIST_MEN(n1707),
    .A_BIST_WEN(n1708),
    .A_BIST_REN(n1709),
    .A_BIST_ADDR(n1710),
    .A_BIST_DIN(n1711),
    .A_BIST_BM(n1712),
    .A_DOUT(\row_n2_inst.A_DOUT ));
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:86:49  */
  assign n1701 = n1665[63:48]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:89:24  */
  assign n1704 = wr_mask[31:16]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:99:60  */
  assign n1714 = n1665[66]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:99:66  */
  assign n1715 = ~n1714;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:99:42  */
  assign n1716 = n1715 ? 8'b00000000 : 8'b11111111;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:100:63  */
  assign n1719 = n1665[67]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:100:71  */
  assign n1720 = ~n1719;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:100:45  */
  assign n1721 = n1720 ? 8'b00000000 : 8'b11111111;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:105:34  */
  assign n1724 = n1665[13:2]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:111:16  */
  assign n1726 = ~rstn_i;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:115:34  */
  assign n1729 = n1665[68]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:115:57  */
  assign n1730 = n1665[69]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:115:43  */
  assign n1731 = ~n1730;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:115:38  */
  assign n1732 = n1729 & n1731;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:116:34  */
  assign n1733 = n1665[68]; // extract
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:120:46  */
  assign n1741 = rden ? rdata : 32'b00000000000000000000000000000000;
  assign n1744 = {\row_n2_inst.A_DOUT , \row_n1_inst.A_DOUT };
  assign n1745 = {n1721, n1716, n1698, n1693};
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:114:5  */
  always @(posedge clk_i or posedge n1726)
    if (n1726)
      n1746 <= 1'b0;
    else
      n1746 <= n1732;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:114:5  */
  always @(posedge clk_i or posedge n1726)
    if (n1726)
      n1748 <= 1'b0;
    else
      n1748 <= n1733;
  /* ../../src/hdl/sg13g2/neorv32_dmem.vhd:111:5  */
  assign n1749 = {1'b0, n1748, n1741};
endmodule

module neorv32_bus_gateway_15_16384_16384_268435456_2097152_d3c572afed0908e1a530126dd188e3360efa598d
  (input  clk_i,
   input  rstn_i,
   input  [31:0] \req_i_req_i[addr] ,
   input  [31:0] \req_i_req_i[data] ,
   input  [3:0] \req_i_req_i[ben] ,
   input  \req_i_req_i[stb] ,
   input  \req_i_req_i[rw] ,
   input  \req_i_req_i[src] ,
   input  \req_i_req_i[priv] ,
   input  \req_i_req_i[amo] ,
   input  [3:0] \req_i_req_i[amoop] ,
   input  \req_i_req_i[fence] ,
   input  \req_i_req_i[sleep] ,
   input  \req_i_req_i[debug] ,
   input  [31:0] \a_rsp_i_a_rsp_i[data] ,
   input  \a_rsp_i_a_rsp_i[ack] ,
   input  \a_rsp_i_a_rsp_i[err] ,
   input  [31:0] \b_rsp_i_b_rsp_i[data] ,
   input  \b_rsp_i_b_rsp_i[ack] ,
   input  \b_rsp_i_b_rsp_i[err] ,
   input  [31:0] \c_rsp_i_c_rsp_i[data] ,
   input  \c_rsp_i_c_rsp_i[ack] ,
   input  \c_rsp_i_c_rsp_i[err] ,
   input  [31:0] \d_rsp_i_d_rsp_i[data] ,
   input  \d_rsp_i_d_rsp_i[ack] ,
   input  \d_rsp_i_d_rsp_i[err] ,
   input  [31:0] \x_rsp_i_x_rsp_i[data] ,
   input  \x_rsp_i_x_rsp_i[ack] ,
   input  \x_rsp_i_x_rsp_i[err] ,
   output [31:0] \rsp_o_rsp_o[data] ,
   output \rsp_o_rsp_o[ack] ,
   output \rsp_o_rsp_o[err] ,
   output [31:0] \a_req_o_a_req_o[addr] ,
   output [31:0] \a_req_o_a_req_o[data] ,
   output [3:0] \a_req_o_a_req_o[ben] ,
   output \a_req_o_a_req_o[stb] ,
   output \a_req_o_a_req_o[rw] ,
   output \a_req_o_a_req_o[src] ,
   output \a_req_o_a_req_o[priv] ,
   output \a_req_o_a_req_o[amo] ,
   output [3:0] \a_req_o_a_req_o[amoop] ,
   output \a_req_o_a_req_o[fence] ,
   output \a_req_o_a_req_o[sleep] ,
   output \a_req_o_a_req_o[debug] ,
   output [31:0] \b_req_o_b_req_o[addr] ,
   output [31:0] \b_req_o_b_req_o[data] ,
   output [3:0] \b_req_o_b_req_o[ben] ,
   output \b_req_o_b_req_o[stb] ,
   output \b_req_o_b_req_o[rw] ,
   output \b_req_o_b_req_o[src] ,
   output \b_req_o_b_req_o[priv] ,
   output \b_req_o_b_req_o[amo] ,
   output [3:0] \b_req_o_b_req_o[amoop] ,
   output \b_req_o_b_req_o[fence] ,
   output \b_req_o_b_req_o[sleep] ,
   output \b_req_o_b_req_o[debug] ,
   output [31:0] \c_req_o_c_req_o[addr] ,
   output [31:0] \c_req_o_c_req_o[data] ,
   output [3:0] \c_req_o_c_req_o[ben] ,
   output \c_req_o_c_req_o[stb] ,
   output \c_req_o_c_req_o[rw] ,
   output \c_req_o_c_req_o[src] ,
   output \c_req_o_c_req_o[priv] ,
   output \c_req_o_c_req_o[amo] ,
   output [3:0] \c_req_o_c_req_o[amoop] ,
   output \c_req_o_c_req_o[fence] ,
   output \c_req_o_c_req_o[sleep] ,
   output \c_req_o_c_req_o[debug] ,
   output [31:0] \d_req_o_d_req_o[addr] ,
   output [31:0] \d_req_o_d_req_o[data] ,
   output [3:0] \d_req_o_d_req_o[ben] ,
   output \d_req_o_d_req_o[stb] ,
   output \d_req_o_d_req_o[rw] ,
   output \d_req_o_d_req_o[src] ,
   output \d_req_o_d_req_o[priv] ,
   output \d_req_o_d_req_o[amo] ,
   output [3:0] \d_req_o_d_req_o[amoop] ,
   output \d_req_o_d_req_o[fence] ,
   output \d_req_o_d_req_o[sleep] ,
   output \d_req_o_d_req_o[debug] ,
   output [31:0] \x_req_o_x_req_o[addr] ,
   output [31:0] \x_req_o_x_req_o[data] ,
   output [3:0] \x_req_o_x_req_o[ben] ,
   output \x_req_o_x_req_o[stb] ,
   output \x_req_o_x_req_o[rw] ,
   output \x_req_o_x_req_o[src] ,
   output \x_req_o_x_req_o[priv] ,
   output \x_req_o_x_req_o[amo] ,
   output [3:0] \x_req_o_x_req_o[amoop] ,
   output \x_req_o_x_req_o[fence] ,
   output \x_req_o_x_req_o[sleep] ,
   output \x_req_o_x_req_o[debug] );
  wire [79:0] n1365;
  wire [31:0] n1367;
  wire n1368;
  wire n1369;
  wire [31:0] n1371;
  wire [31:0] n1372;
  wire [3:0] n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire [3:0] n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire [33:0] n1383;
  wire [31:0] n1385;
  wire [31:0] n1386;
  wire [3:0] n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire [3:0] n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire [33:0] n1397;
  wire [31:0] n1399;
  wire [31:0] n1400;
  wire [3:0] n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire [3:0] n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire [33:0] n1411;
  wire [31:0] n1413;
  wire [31:0] n1414;
  wire [3:0] n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire [3:0] n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire [33:0] n1425;
  wire [31:0] n1427;
  wire [31:0] n1428;
  wire [3:0] n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire [3:0] n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire [33:0] n1439;
  wire [4:0] port_sel;
  wire [399:0] port_req;
  wire [169:0] port_rsp;
  wire [33:0] int_rsp;
  wire [7:0] keeper;
  wire n1442;
  wire [17:0] n1446;
  wire n1449;
  wire n1451;
  wire n1452;
  wire [3:0] n1456;
  wire n1459;
  wire n1461;
  wire n1462;
  wire [10:0] n1466;
  wire n1469;
  wire n1471;
  wire n1472;
  wire [3:0] n1475;
  wire n1477;
  wire n1479;
  wire n1480;
  wire [79:0] n1482;
  wire [79:0] n1483;
  wire [79:0] n1484;
  wire [79:0] n1485;
  wire [79:0] n1486;
  wire n1489;
  wire n1490;
  wire n1491;
  wire [10:0] n1492;
  wire [67:0] n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire [10:0] n1497;
  wire [67:0] n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire [10:0] n1502;
  wire [67:0] n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire [10:0] n1507;
  wire [67:0] n1508;
  localparam [33:0] n1512 = 34'b0000000000000000000000000000000000;
  wire [31:0] n1513;
  wire [31:0] n1515;
  wire [31:0] n1516;
  localparam [33:0] n1517 = 34'b0000000000000000000000000000000000;
  wire [1:0] n1518;
  wire [33:0] n1519;
  wire n1520;
  wire n1522;
  wire n1523;
  wire n1524;
  wire [33:0] n1525;
  wire n1526;
  wire n1528;
  wire n1529;
  wire [33:0] n1530;
  wire [31:0] n1531;
  wire [31:0] n1533;
  wire [31:0] n1534;
  wire [33:0] n1535;
  wire n1536;
  wire n1538;
  wire n1539;
  wire [33:0] n1540;
  wire n1541;
  wire n1543;
  wire n1544;
  wire [33:0] n1545;
  wire [31:0] n1546;
  wire [31:0] n1548;
  wire [31:0] n1549;
  wire [33:0] n1550;
  wire n1551;
  wire n1553;
  wire n1554;
  wire [33:0] n1555;
  wire n1556;
  wire n1558;
  wire n1559;
  wire [33:0] n1560;
  wire [31:0] n1561;
  wire [31:0] n1563;
  wire [31:0] n1564;
  wire [33:0] n1565;
  wire n1566;
  wire n1568;
  wire n1569;
  wire [33:0] n1570;
  wire n1571;
  wire n1573;
  wire n1574;
  wire [33:0] n1575;
  wire [31:0] n1578;
  wire n1579;
  wire n1580;
  wire n1582;
  wire [4:0] n1591;
  wire n1597;
  wire n1599;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1612;
  wire [4:0] n1613;
  wire [4:0] n1615;
  wire n1616;
  wire n1624;
  wire n1626;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1643;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire [6:0] n1649;
  wire [5:0] n1650;
  wire [5:0] n1651;
  wire [5:0] n1652;
  wire n1653;
  wire n1654;
  wire [7:0] n1655;
  wire [7:0] n1657;
  wire [4:0] n1660;
  wire [399:0] n1661;
  wire [169:0] n1662;
  reg [7:0] n1663;
  wire [33:0] n1664;
  assign \rsp_o_rsp_o[data]  = n1367; //(module output)
  assign \rsp_o_rsp_o[ack]  = n1368; //(module output)
  assign \rsp_o_rsp_o[err]  = n1369; //(module output)
  assign \a_req_o_a_req_o[addr]  = n1371; //(module output)
  assign \a_req_o_a_req_o[data]  = n1372; //(module output)
  assign \a_req_o_a_req_o[ben]  = n1373; //(module output)
  assign \a_req_o_a_req_o[stb]  = n1374; //(module output)
  assign \a_req_o_a_req_o[rw]  = n1375; //(module output)
  assign \a_req_o_a_req_o[src]  = n1376; //(module output)
  assign \a_req_o_a_req_o[priv]  = n1377; //(module output)
  assign \a_req_o_a_req_o[amo]  = n1378; //(module output)
  assign \a_req_o_a_req_o[amoop]  = n1379; //(module output)
  assign \a_req_o_a_req_o[fence]  = n1380; //(module output)
  assign \a_req_o_a_req_o[sleep]  = n1381; //(module output)
  assign \a_req_o_a_req_o[debug]  = n1382; //(module output)
  assign \b_req_o_b_req_o[addr]  = n1385; //(module output)
  assign \b_req_o_b_req_o[data]  = n1386; //(module output)
  assign \b_req_o_b_req_o[ben]  = n1387; //(module output)
  assign \b_req_o_b_req_o[stb]  = n1388; //(module output)
  assign \b_req_o_b_req_o[rw]  = n1389; //(module output)
  assign \b_req_o_b_req_o[src]  = n1390; //(module output)
  assign \b_req_o_b_req_o[priv]  = n1391; //(module output)
  assign \b_req_o_b_req_o[amo]  = n1392; //(module output)
  assign \b_req_o_b_req_o[amoop]  = n1393; //(module output)
  assign \b_req_o_b_req_o[fence]  = n1394; //(module output)
  assign \b_req_o_b_req_o[sleep]  = n1395; //(module output)
  assign \b_req_o_b_req_o[debug]  = n1396; //(module output)
  assign \c_req_o_c_req_o[addr]  = n1399; //(module output)
  assign \c_req_o_c_req_o[data]  = n1400; //(module output)
  assign \c_req_o_c_req_o[ben]  = n1401; //(module output)
  assign \c_req_o_c_req_o[stb]  = n1402; //(module output)
  assign \c_req_o_c_req_o[rw]  = n1403; //(module output)
  assign \c_req_o_c_req_o[src]  = n1404; //(module output)
  assign \c_req_o_c_req_o[priv]  = n1405; //(module output)
  assign \c_req_o_c_req_o[amo]  = n1406; //(module output)
  assign \c_req_o_c_req_o[amoop]  = n1407; //(module output)
  assign \c_req_o_c_req_o[fence]  = n1408; //(module output)
  assign \c_req_o_c_req_o[sleep]  = n1409; //(module output)
  assign \c_req_o_c_req_o[debug]  = n1410; //(module output)
  assign \d_req_o_d_req_o[addr]  = n1413; //(module output)
  assign \d_req_o_d_req_o[data]  = n1414; //(module output)
  assign \d_req_o_d_req_o[ben]  = n1415; //(module output)
  assign \d_req_o_d_req_o[stb]  = n1416; //(module output)
  assign \d_req_o_d_req_o[rw]  = n1417; //(module output)
  assign \d_req_o_d_req_o[src]  = n1418; //(module output)
  assign \d_req_o_d_req_o[priv]  = n1419; //(module output)
  assign \d_req_o_d_req_o[amo]  = n1420; //(module output)
  assign \d_req_o_d_req_o[amoop]  = n1421; //(module output)
  assign \d_req_o_d_req_o[fence]  = n1422; //(module output)
  assign \d_req_o_d_req_o[sleep]  = n1423; //(module output)
  assign \d_req_o_d_req_o[debug]  = n1424; //(module output)
  assign \x_req_o_x_req_o[addr]  = n1427; //(module output)
  assign \x_req_o_x_req_o[data]  = n1428; //(module output)
  assign \x_req_o_x_req_o[ben]  = n1429; //(module output)
  assign \x_req_o_x_req_o[stb]  = n1430; //(module output)
  assign \x_req_o_x_req_o[rw]  = n1431; //(module output)
  assign \x_req_o_x_req_o[src]  = n1432; //(module output)
  assign \x_req_o_x_req_o[priv]  = n1433; //(module output)
  assign \x_req_o_x_req_o[amo]  = n1434; //(module output)
  assign \x_req_o_x_req_o[amoop]  = n1435; //(module output)
  assign \x_req_o_x_req_o[fence]  = n1436; //(module output)
  assign \x_req_o_x_req_o[sleep]  = n1437; //(module output)
  assign \x_req_o_x_req_o[debug]  = n1438; //(module output)
  assign n1365 = {\req_i_req_i[debug] , \req_i_req_i[sleep] , \req_i_req_i[fence] , \req_i_req_i[amoop] , \req_i_req_i[amo] , \req_i_req_i[priv] , \req_i_req_i[src] , \req_i_req_i[rw] , \req_i_req_i[stb] , \req_i_req_i[ben] , \req_i_req_i[data] , \req_i_req_i[addr] };
  assign n1367 = n1664[31:0]; // extract
  assign n1368 = n1664[32]; // extract
  assign n1369 = n1664[33]; // extract
  assign n1371 = n1482[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:48:3  */
  assign n1372 = n1482[63:32]; // extract
  assign n1373 = n1482[67:64]; // extract
  assign n1374 = n1482[68]; // extract
  assign n1375 = n1482[69]; // extract
  assign n1376 = n1482[70]; // extract
  assign n1377 = n1482[71]; // extract
  assign n1378 = n1482[72]; // extract
  assign n1379 = n1482[76:73]; // extract
  assign n1380 = n1482[77]; // extract
  assign n1381 = n1482[78]; // extract
  assign n1382 = n1482[79]; // extract
  assign n1383 = {\a_rsp_i_a_rsp_i[err] , \a_rsp_i_a_rsp_i[ack] , \a_rsp_i_a_rsp_i[data] };
  assign n1385 = n1483[31:0]; // extract
  assign n1386 = n1483[63:32]; // extract
  assign n1387 = n1483[67:64]; // extract
  assign n1388 = n1483[68]; // extract
  assign n1389 = n1483[69]; // extract
  assign n1390 = n1483[70]; // extract
  assign n1391 = n1483[71]; // extract
  assign n1392 = n1483[72]; // extract
  assign n1393 = n1483[76:73]; // extract
  assign n1394 = n1483[77]; // extract
  assign n1395 = n1483[78]; // extract
  assign n1396 = n1483[79]; // extract
  assign n1397 = {\b_rsp_i_b_rsp_i[err] , \b_rsp_i_b_rsp_i[ack] , \b_rsp_i_b_rsp_i[data] };
  assign n1399 = n1484[31:0]; // extract
  assign n1400 = n1484[63:32]; // extract
  assign n1401 = n1484[67:64]; // extract
  assign n1402 = n1484[68]; // extract
  assign n1403 = n1484[69]; // extract
  assign n1404 = n1484[70]; // extract
  assign n1405 = n1484[71]; // extract
  assign n1406 = n1484[72]; // extract
  assign n1407 = n1484[76:73]; // extract
  assign n1408 = n1484[77]; // extract
  assign n1409 = n1484[78]; // extract
  assign n1410 = n1484[79]; // extract
  assign n1411 = {\c_rsp_i_c_rsp_i[err] , \c_rsp_i_c_rsp_i[ack] , \c_rsp_i_c_rsp_i[data] };
  assign n1413 = n1485[31:0]; // extract
  assign n1414 = n1485[63:32]; // extract
  assign n1415 = n1485[67:64]; // extract
  assign n1416 = n1485[68]; // extract
  assign n1417 = n1485[69]; // extract
  assign n1418 = n1485[70]; // extract
  assign n1419 = n1485[71]; // extract
  assign n1420 = n1485[72]; // extract
  assign n1421 = n1485[76:73]; // extract
  assign n1422 = n1485[77]; // extract
  assign n1423 = n1485[78]; // extract
  assign n1424 = n1485[79]; // extract
  assign n1425 = {\d_rsp_i_d_rsp_i[err] , \d_rsp_i_d_rsp_i[ack] , \d_rsp_i_d_rsp_i[data] };
  assign n1427 = n1486[31:0]; // extract
  assign n1428 = n1486[63:32]; // extract
  assign n1429 = n1486[67:64]; // extract
  assign n1430 = n1486[68]; // extract
  assign n1431 = n1486[69]; // extract
  assign n1432 = n1486[70]; // extract
  assign n1433 = n1486[71]; // extract
  assign n1434 = n1486[72]; // extract
  assign n1435 = n1486[76:73]; // extract
  assign n1436 = n1486[77]; // extract
  assign n1437 = n1486[78]; // extract
  assign n1438 = n1486[79]; // extract
  assign n1439 = {\x_rsp_i_x_rsp_i[err] , \x_rsp_i_x_rsp_i[ack] , \x_rsp_i_x_rsp_i[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:367:10  */
  assign port_sel = n1660; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:381:10  */
  assign port_req = n1661; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:382:10  */
  assign port_rsp = n1662; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:385:10  */
  assign int_rsp = n1575; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:394:10  */
  assign keeper = n1663; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:400:22  */
  assign n1442 = 1'b0 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:401:51  */
  assign n1446 = n1365[31:14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:401:84  */
  assign n1449 = n1446 == 18'b100000000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:401:36  */
  assign n1451 = n1449 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:401:22  */
  assign n1452 = n1451 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:402:51  */
  assign n1456 = n1365[31:28]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:402:84  */
  assign n1459 = n1456 == 4'b1110;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:402:36  */
  assign n1461 = n1459 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:402:22  */
  assign n1462 = n1461 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:403:51  */
  assign n1466 = n1365[31:21]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:403:84  */
  assign n1469 = n1466 == 11'b11111111111;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:403:36  */
  assign n1471 = n1469 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:403:22  */
  assign n1472 = n1471 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:406:49  */
  assign n1475 = port_sel[3:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:406:62  */
  assign n1477 = n1475 == 4'b0000;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:406:36  */
  assign n1479 = n1477 & 1'b1;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:406:22  */
  assign n1480 = n1479 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:411:22  */
  assign n1482 = port_req[399:320]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:412:22  */
  assign n1483 = port_req[319:240]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:413:22  */
  assign n1484 = port_req[239:160]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:414:22  */
  assign n1485 = port_req[159:80]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:415:22  */
  assign n1486 = port_req[79:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:36  */
  assign n1489 = port_sel[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:50  */
  assign n1490 = n1365[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:40  */
  assign n1491 = n1489 & n1490;
  assign n1492 = n1365[79:69]; // extract
  assign n1493 = n1365[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:36  */
  assign n1494 = port_sel[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:50  */
  assign n1495 = n1365[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:40  */
  assign n1496 = n1494 & n1495;
  assign n1497 = n1365[79:69]; // extract
  assign n1498 = n1365[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:36  */
  assign n1499 = port_sel[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:50  */
  assign n1500 = n1365[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:40  */
  assign n1501 = n1499 & n1500;
  assign n1502 = n1365[79:69]; // extract
  assign n1503 = n1365[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:36  */
  assign n1504 = port_sel[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:50  */
  assign n1505 = n1365[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:424:40  */
  assign n1506 = n1504 & n1505;
  assign n1507 = n1365[79:69]; // extract
  assign n1508 = n1365[67:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:29  */
  assign n1513 = n1512[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:49  */
  assign n1515 = port_rsp[133:102]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:34  */
  assign n1516 = n1513 | n1515;
  assign n1518 = n1517[33:32]; // extract
  assign n1519 = {n1518, n1516};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:29  */
  assign n1520 = n1519[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:49  */
  assign n1522 = port_rsp[134]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:34  */
  assign n1523 = n1520 | n1522;
  assign n1524 = n1517[33]; // extract
  assign n1525 = {n1524, n1523, n1516};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:29  */
  assign n1526 = n1525[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:49  */
  assign n1528 = port_rsp[135]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:34  */
  assign n1529 = n1526 | n1528;
  assign n1530 = {n1529, n1523, n1516};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:29  */
  assign n1531 = n1530[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:49  */
  assign n1533 = port_rsp[99:68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:34  */
  assign n1534 = n1531 | n1533;
  assign n1535 = {n1529, n1523, n1534};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:29  */
  assign n1536 = n1535[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:49  */
  assign n1538 = port_rsp[100]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:34  */
  assign n1539 = n1536 | n1538;
  assign n1540 = {n1529, n1539, n1534};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:29  */
  assign n1541 = n1540[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:49  */
  assign n1543 = port_rsp[101]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:34  */
  assign n1544 = n1541 | n1543;
  assign n1545 = {n1544, n1539, n1534};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:29  */
  assign n1546 = n1545[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:49  */
  assign n1548 = port_rsp[65:34]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:34  */
  assign n1549 = n1546 | n1548;
  assign n1550 = {n1544, n1539, n1549};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:29  */
  assign n1551 = n1550[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:49  */
  assign n1553 = port_rsp[66]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:34  */
  assign n1554 = n1551 | n1553;
  assign n1555 = {n1544, n1554, n1549};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:29  */
  assign n1556 = n1555[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:49  */
  assign n1558 = port_rsp[67]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:34  */
  assign n1559 = n1556 | n1558;
  assign n1560 = {n1559, n1554, n1549};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:29  */
  assign n1561 = n1560[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:49  */
  assign n1563 = port_rsp[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:436:34  */
  assign n1564 = n1561 | n1563;
  assign n1565 = {n1559, n1554, n1564};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:29  */
  assign n1566 = n1565[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:49  */
  assign n1568 = port_rsp[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:437:34  */
  assign n1569 = n1566 | n1568;
  assign n1570 = {n1559, n1569, n1564};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:29  */
  assign n1571 = n1570[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:49  */
  assign n1573 = port_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:438:34  */
  assign n1574 = n1571 | n1573;
  assign n1575 = {n1574, n1569, n1564};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:445:25  */
  assign n1578 = int_rsp[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:446:25  */
  assign n1579 = int_rsp[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:447:24  */
  assign n1580 = keeper[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:454:16  */
  assign n1582 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:461:43  */
  assign n1591 = port_sel & 5'b10100;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1597 = n1591[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1599 = 1'b0 | n1597;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1601 = n1591[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1602 = n1599 | n1601;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1603 = n1591[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1604 = n1602 | n1603;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1605 = n1591[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1606 = n1604 | n1605;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1607 = n1591[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1608 = n1606 | n1607;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:462:18  */
  assign n1609 = keeper[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:462:23  */
  assign n1610 = ~n1609;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:464:30  */
  assign n1612 = n1365[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:466:57  */
  assign n1613 = keeper[5:1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:466:62  */
  assign n1615 = n1613 - 5'b00001;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:467:21  */
  assign n1616 = int_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1624 = keeper[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1626 = 1'b0 | n1624;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1628 = keeper[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1629 = n1626 | n1628;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1630 = keeper[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1631 = n1629 | n1630;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1632 = keeper[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1633 = n1631 | n1632;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n1634 = keeper[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n1635 = n1633 | n1634;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:467:61  */
  assign n1636 = ~n1635;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:467:80  */
  assign n1637 = keeper[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:467:85  */
  assign n1638 = ~n1637;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:467:68  */
  assign n1639 = n1638 & n1636;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:467:32  */
  assign n1640 = n1616 | n1639;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:470:24  */
  assign n1643 = int_rsp[32]; // extract
  assign n1645 = keeper[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:470:9  */
  assign n1646 = n1643 ? 1'b0 : n1645;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:467:9  */
  assign n1647 = n1640 ? 1'b0 : n1646;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:467:9  */
  assign n1648 = n1640 ? 1'b1 : 1'b0;
  assign n1649 = {n1648, n1615, n1647};
  assign n1650 = {5'b01111, n1612};
  assign n1651 = n1649[5:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:462:7  */
  assign n1652 = n1610 ? n1650 : n1651;
  assign n1653 = n1649[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:462:7  */
  assign n1654 = n1610 ? 1'b0 : n1653;
  assign n1655 = {n1608, n1654, n1652};
  assign n1657 = {1'b0, 1'b0, 5'b00000, 1'b0};
  assign n1660 = {n1480, n1472, n1462, n1452, n1442};
  assign n1661 = {80'b01000000000000000000000000000000000000000000000000000000000000000000000000000000, n1492, n1491, n1493, n1497, n1496, n1498, n1502, n1501, n1503, n1507, n1506, n1508};
  assign n1662 = {n1383, n1397, n1411, n1425, n1439};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:459:5  */
  always @(posedge clk_i or posedge n1582)
    if (n1582)
      n1663 <= n1657;
    else
      n1663 <= n1655;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:454:5  */
  assign n1664 = {n1580, n1579, n1578};
endmodule

module neorv32_bus_switch_2547cc736e951fa4919853c43ae890861a3b3264
  (input  clk_i,
   input  rstn_i,
   input  a_lock_i,
   input  [31:0] \a_req_i_a_req_i[addr] ,
   input  [31:0] \a_req_i_a_req_i[data] ,
   input  [3:0] \a_req_i_a_req_i[ben] ,
   input  \a_req_i_a_req_i[stb] ,
   input  \a_req_i_a_req_i[rw] ,
   input  \a_req_i_a_req_i[src] ,
   input  \a_req_i_a_req_i[priv] ,
   input  \a_req_i_a_req_i[amo] ,
   input  [3:0] \a_req_i_a_req_i[amoop] ,
   input  \a_req_i_a_req_i[fence] ,
   input  \a_req_i_a_req_i[sleep] ,
   input  \a_req_i_a_req_i[debug] ,
   input  [31:0] \b_req_i_b_req_i[addr] ,
   input  [31:0] \b_req_i_b_req_i[data] ,
   input  [3:0] \b_req_i_b_req_i[ben] ,
   input  \b_req_i_b_req_i[stb] ,
   input  \b_req_i_b_req_i[rw] ,
   input  \b_req_i_b_req_i[src] ,
   input  \b_req_i_b_req_i[priv] ,
   input  \b_req_i_b_req_i[amo] ,
   input  [3:0] \b_req_i_b_req_i[amoop] ,
   input  \b_req_i_b_req_i[fence] ,
   input  \b_req_i_b_req_i[sleep] ,
   input  \b_req_i_b_req_i[debug] ,
   input  [31:0] \x_rsp_i_x_rsp_i[data] ,
   input  \x_rsp_i_x_rsp_i[ack] ,
   input  \x_rsp_i_x_rsp_i[err] ,
   output [31:0] \a_rsp_o_a_rsp_o[data] ,
   output \a_rsp_o_a_rsp_o[ack] ,
   output \a_rsp_o_a_rsp_o[err] ,
   output [31:0] \b_rsp_o_b_rsp_o[data] ,
   output \b_rsp_o_b_rsp_o[ack] ,
   output \b_rsp_o_b_rsp_o[err] ,
   output [31:0] \x_req_o_x_req_o[addr] ,
   output [31:0] \x_req_o_x_req_o[data] ,
   output [3:0] \x_req_o_x_req_o[ben] ,
   output \x_req_o_x_req_o[stb] ,
   output \x_req_o_x_req_o[rw] ,
   output \x_req_o_x_req_o[src] ,
   output \x_req_o_x_req_o[priv] ,
   output \x_req_o_x_req_o[amo] ,
   output [3:0] \x_req_o_x_req_o[amoop] ,
   output \x_req_o_x_req_o[fence] ,
   output \x_req_o_x_req_o[sleep] ,
   output \x_req_o_x_req_o[debug] );
  wire [79:0] n1195;
  wire [31:0] n1197;
  wire n1198;
  wire n1199;
  wire [79:0] n1200;
  wire [31:0] n1202;
  wire n1203;
  wire n1204;
  wire [31:0] n1206;
  wire [31:0] n1207;
  wire [3:0] n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire [3:0] n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire [33:0] n1218;
  wire [1:0] state;
  wire [1:0] state_nxt;
  wire a_req;
  wire b_req;
  wire sel;
  wire stb;
  wire n1220;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1227;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1233;
  wire n1245;
  wire n1246;
  wire n1247;
  wire [1:0] n1249;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire [1:0] n1256;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire [1:0] n1266;
  wire n1269;
  wire n1272;
  wire [1:0] n1274;
  wire n1276;
  wire n1278;
  wire [1:0] n1279;
  reg [1:0] n1280;
  reg n1283;
  reg n1286;
  wire [31:0] n1289;
  wire n1290;
  wire [31:0] n1291;
  wire [31:0] n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire [3:0] n1297;
  wire n1298;
  wire [3:0] n1299;
  wire [3:0] n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire [31:0] n1323;
  wire [31:0] n1325;
  wire [31:0] n1326;
  wire [31:0] n1328;
  wire [31:0] n1329;
  wire n1330;
  wire [31:0] n1331;
  wire [31:0] n1332;
  wire [3:0] n1333;
  wire [3:0] n1335;
  wire [3:0] n1336;
  wire [3:0] n1338;
  wire [3:0] n1339;
  wire n1340;
  wire [3:0] n1341;
  wire [3:0] n1342;
  wire [31:0] n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1348;
  wire n1349;
  wire n1350;
  wire [31:0] n1352;
  wire n1353;
  wire n1354;
  wire n1356;
  wire n1357;
  reg [1:0] n1359;
  reg n1360;
  reg n1361;
  wire [33:0] n1362;
  wire [33:0] n1363;
  wire [79:0] n1364;
  assign \a_rsp_o_a_rsp_o[data]  = n1197; //(module output)
  assign \a_rsp_o_a_rsp_o[ack]  = n1198; //(module output)
  assign \a_rsp_o_a_rsp_o[err]  = n1199; //(module output)
  assign \b_rsp_o_b_rsp_o[data]  = n1202; //(module output)
  assign \b_rsp_o_b_rsp_o[ack]  = n1203; //(module output)
  assign \b_rsp_o_b_rsp_o[err]  = n1204; //(module output)
  assign \x_req_o_x_req_o[addr]  = n1206; //(module output)
  assign \x_req_o_x_req_o[data]  = n1207; //(module output)
  assign \x_req_o_x_req_o[ben]  = n1208; //(module output)
  assign \x_req_o_x_req_o[stb]  = n1209; //(module output)
  assign \x_req_o_x_req_o[rw]  = n1210; //(module output)
  assign \x_req_o_x_req_o[src]  = n1211; //(module output)
  assign \x_req_o_x_req_o[priv]  = n1212; //(module output)
  assign \x_req_o_x_req_o[amo]  = n1213; //(module output)
  assign \x_req_o_x_req_o[amoop]  = n1214; //(module output)
  assign \x_req_o_x_req_o[fence]  = n1215; //(module output)
  assign \x_req_o_x_req_o[sleep]  = n1216; //(module output)
  assign \x_req_o_x_req_o[debug]  = n1217; //(module output)
  assign n1195 = {\a_req_i_a_req_i[debug] , \a_req_i_a_req_i[sleep] , \a_req_i_a_req_i[fence] , \a_req_i_a_req_i[amoop] , \a_req_i_a_req_i[amo] , \a_req_i_a_req_i[priv] , \a_req_i_a_req_i[src] , \a_req_i_a_req_i[rw] , \a_req_i_a_req_i[stb] , \a_req_i_a_req_i[ben] , \a_req_i_a_req_i[data] , \a_req_i_a_req_i[addr] };
  assign n1197 = n1362[31:0]; // extract
  assign n1198 = n1362[32]; // extract
  assign n1199 = n1362[33]; // extract
  assign n1200 = {\b_req_i_b_req_i[debug] , \b_req_i_b_req_i[sleep] , \b_req_i_b_req_i[fence] , \b_req_i_b_req_i[amoop] , \b_req_i_b_req_i[amo] , \b_req_i_b_req_i[priv] , \b_req_i_b_req_i[src] , \b_req_i_b_req_i[rw] , \b_req_i_b_req_i[stb] , \b_req_i_b_req_i[ben] , \b_req_i_b_req_i[data] , \b_req_i_b_req_i[addr] };
  assign n1202 = n1363[31:0]; // extract
  assign n1203 = n1363[32]; // extract
  assign n1204 = n1363[33]; // extract
  assign n1206 = n1364[31:0]; // extract
  assign n1207 = n1364[63:32]; // extract
  assign n1208 = n1364[67:64]; // extract
  assign n1209 = n1364[68]; // extract
  assign n1210 = n1364[69]; // extract
  assign n1211 = n1364[70]; // extract
  assign n1212 = n1364[71]; // extract
  assign n1213 = n1364[72]; // extract
  assign n1214 = n1364[76:73]; // extract
  assign n1215 = n1364[77]; // extract
  assign n1216 = n1364[78]; // extract
  assign n1217 = n1364[79]; // extract
  assign n1218 = {\x_rsp_i_x_rsp_i[err] , \x_rsp_i_x_rsp_i[ack] , \x_rsp_i_x_rsp_i[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:40:10  */
  assign state = n1359; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:40:17  */
  assign state_nxt = n1280; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:41:10  */
  assign a_req = n1360; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:41:17  */
  assign b_req = n1361; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:42:10  */
  assign sel = n1283; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:42:17  */
  assign stb = n1286; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:50:16  */
  assign n1220 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:56:17  */
  assign n1223 = state == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:59:35  */
  assign n1224 = n1195[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:59:24  */
  assign n1225 = a_req | n1224;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:56:7  */
  assign n1227 = n1223 ? 1'b0 : n1225;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:61:17  */
  assign n1229 = state == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:64:35  */
  assign n1230 = n1200[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:64:24  */
  assign n1231 = b_req | n1230;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:61:7  */
  assign n1233 = n1229 ? 1'b0 : n1231;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:87:23  */
  assign n1245 = n1218[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:87:46  */
  assign n1246 = n1218[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:87:34  */
  assign n1247 = n1245 | n1246;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:87:11  */
  assign n1249 = n1247 ? 2'b00 : state;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:84:9  */
  assign n1251 = state == 2'b01;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:94:23  */
  assign n1252 = n1218[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:94:46  */
  assign n1253 = n1218[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:94:34  */
  assign n1254 = n1252 | n1253;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:94:11  */
  assign n1256 = n1254 ? 2'b00 : state;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:91:9  */
  assign n1258 = state == 2'b11;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:100:23  */
  assign n1259 = n1195[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:100:34  */
  assign n1260 = n1259 | a_req;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:104:27  */
  assign n1261 = n1200[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:104:38  */
  assign n1262 = n1261 | b_req;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:104:70  */
  assign n1263 = ~a_lock_i;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:104:56  */
  assign n1264 = n1263 & n1262;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:104:11  */
  assign n1266 = n1264 ? 2'b11 : state;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:104:11  */
  assign n1269 = n1264 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:104:11  */
  assign n1272 = n1264 ? 1'b1 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:100:11  */
  assign n1274 = n1260 ? 2'b01 : n1266;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:100:11  */
  assign n1276 = n1260 ? 1'b0 : n1269;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:100:11  */
  assign n1278 = n1260 ? 1'b1 : n1272;
  assign n1279 = {n1258, n1251};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:82:7  */
  always @*
    case (n1279)
      2'b10: n1280 = n1256;
      2'b01: n1280 = n1249;
      default: n1280 = n1274;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:82:7  */
  always @*
    case (n1279)
      2'b10: n1283 = 1'b1;
      2'b01: n1283 = 1'b0;
      default: n1283 = n1276;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:82:7  */
  always @*
    case (n1279)
      2'b10: n1286 = 1'b0;
      2'b01: n1286 = 1'b0;
      default: n1286 = n1278;
    endcase
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:174:28  */
  assign n1289 = n1195[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:174:44  */
  assign n1290 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:174:34  */
  assign n1291 = n1290 ? n1289 : n1292;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:174:64  */
  assign n1292 = n1200[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:175:28  */
  assign n1293 = n1195[72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:175:44  */
  assign n1294 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:175:34  */
  assign n1295 = n1294 ? n1293 : n1296;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:175:64  */
  assign n1296 = n1200[72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:176:28  */
  assign n1297 = n1195[76:73]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:176:44  */
  assign n1298 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:176:34  */
  assign n1299 = n1298 ? n1297 : n1300;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:176:64  */
  assign n1300 = n1200[76:73]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:177:28  */
  assign n1301 = n1195[71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:177:44  */
  assign n1302 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:177:34  */
  assign n1303 = n1302 ? n1301 : n1304;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:177:64  */
  assign n1304 = n1200[71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:178:28  */
  assign n1305 = n1195[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:178:44  */
  assign n1306 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:178:34  */
  assign n1307 = n1306 ? n1305 : n1308;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:178:64  */
  assign n1308 = n1200[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:179:28  */
  assign n1309 = n1195[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:179:44  */
  assign n1310 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:179:34  */
  assign n1311 = n1310 ? n1309 : n1312;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:179:64  */
  assign n1312 = n1200[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:180:28  */
  assign n1313 = n1195[77]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:180:46  */
  assign n1314 = n1200[77]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:180:34  */
  assign n1315 = n1313 | n1314;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:181:28  */
  assign n1316 = n1195[78]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:181:46  */
  assign n1317 = n1200[78]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:181:34  */
  assign n1318 = n1316 & n1317;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:182:28  */
  assign n1319 = n1195[79]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:182:44  */
  assign n1320 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:182:34  */
  assign n1321 = n1320 ? n1319 : n1322;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:182:64  */
  assign n1322 = n1200[79]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:184:28  */
  assign n1323 = n1200[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:184:34  */
  assign n1325 = 1'b0 ? n1323 : n1328;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:185:28  */
  assign n1326 = n1195[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:184:59  */
  assign n1328 = 1'b1 ? n1326 : n1331;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:186:28  */
  assign n1329 = n1195[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:186:44  */
  assign n1330 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:185:59  */
  assign n1331 = n1330 ? n1329 : n1332;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:186:64  */
  assign n1332 = n1200[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:188:28  */
  assign n1333 = n1200[67:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:188:34  */
  assign n1335 = 1'b0 ? n1333 : n1338;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:189:28  */
  assign n1336 = n1195[67:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:188:59  */
  assign n1338 = 1'b1 ? n1336 : n1341;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:190:28  */
  assign n1339 = n1195[67:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:190:44  */
  assign n1340 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:189:59  */
  assign n1341 = n1340 ? n1339 : n1342;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:190:64  */
  assign n1342 = n1200[67:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:197:27  */
  assign n1343 = n1218[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:198:27  */
  assign n1344 = n1218[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:198:41  */
  assign n1345 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:198:31  */
  assign n1346 = n1345 ? n1344 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:199:27  */
  assign n1348 = n1218[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:199:41  */
  assign n1349 = ~sel;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:199:31  */
  assign n1350 = n1349 ? n1348 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:201:27  */
  assign n1352 = n1218[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:202:27  */
  assign n1353 = n1218[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:202:31  */
  assign n1354 = sel ? n1353 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:203:27  */
  assign n1356 = n1218[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:203:31  */
  assign n1357 = sel ? n1356 : 1'b0;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:54:5  */
  always @(posedge clk_i or posedge n1220)
    if (n1220)
      n1359 <= 2'b00;
    else
      n1359 <= state_nxt;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:54:5  */
  always @(posedge clk_i or posedge n1220)
    if (n1220)
      n1360 <= 1'b0;
    else
      n1360 <= n1227;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:54:5  */
  always @(posedge clk_i or posedge n1220)
    if (n1220)
      n1361 <= 1'b0;
    else
      n1361 <= n1233;
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:50:5  */
  assign n1362 = {n1350, n1346, n1343};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:50:5  */
  assign n1363 = {n1357, n1354, n1352};
  /* ../../ext/neorv32/rtl/core/neorv32_bus.vhd:50:5  */
  assign n1364 = {n1321, n1318, n1315, n1299, n1295, n1303, n1307, n1311, stb, n1335, n1325, n1291};
endmodule

module neorv32_cpu_0_0_4_1_40_f23860951627a2ed8cecb4a83038f47ead6bd96c
  (input  clk_i,
   input  rstn_i,
   input  msi_i,
   input  mei_i,
   input  mti_i,
   input  [15:0] firq_i,
   input  dbi_i,
   input  \icc_rx_i_icc_rx_i[rdy] ,
   input  \icc_rx_i_icc_rx_i[ack] ,
   input  [31:0] \icc_rx_i_icc_rx_i[dat] ,
   input  [31:0] \ibus_rsp_i_ibus_rsp_i[data] ,
   input  \ibus_rsp_i_ibus_rsp_i[ack] ,
   input  \ibus_rsp_i_ibus_rsp_i[err] ,
   input  [31:0] \dbus_rsp_i_dbus_rsp_i[data] ,
   input  \dbus_rsp_i_dbus_rsp_i[ack] ,
   input  \dbus_rsp_i_dbus_rsp_i[err] ,
   output \icc_tx_o_icc_tx_o[rdy] ,
   output \icc_tx_o_icc_tx_o[ack] ,
   output [31:0] \icc_tx_o_icc_tx_o[dat] ,
   output [31:0] \ibus_req_o_ibus_req_o[addr] ,
   output [31:0] \ibus_req_o_ibus_req_o[data] ,
   output [3:0] \ibus_req_o_ibus_req_o[ben] ,
   output \ibus_req_o_ibus_req_o[stb] ,
   output \ibus_req_o_ibus_req_o[rw] ,
   output \ibus_req_o_ibus_req_o[src] ,
   output \ibus_req_o_ibus_req_o[priv] ,
   output \ibus_req_o_ibus_req_o[amo] ,
   output [3:0] \ibus_req_o_ibus_req_o[amoop] ,
   output \ibus_req_o_ibus_req_o[fence] ,
   output \ibus_req_o_ibus_req_o[sleep] ,
   output \ibus_req_o_ibus_req_o[debug] ,
   output [31:0] \dbus_req_o_dbus_req_o[addr] ,
   output [31:0] \dbus_req_o_dbus_req_o[data] ,
   output [3:0] \dbus_req_o_dbus_req_o[ben] ,
   output \dbus_req_o_dbus_req_o[stb] ,
   output \dbus_req_o_dbus_req_o[rw] ,
   output \dbus_req_o_dbus_req_o[src] ,
   output \dbus_req_o_dbus_req_o[priv] ,
   output \dbus_req_o_dbus_req_o[amo] ,
   output [3:0] \dbus_req_o_dbus_req_o[amoop] ,
   output \dbus_req_o_dbus_req_o[fence] ,
   output \dbus_req_o_dbus_req_o[sleep] ,
   output \dbus_req_o_dbus_req_o[debug] );
  wire n1005;
  wire n1006;
  wire [31:0] n1007;
  wire [31:0] n1010;
  wire [31:0] n1011;
  wire [3:0] n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire [3:0] n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire [33:0] n1022;
  wire [31:0] n1024;
  wire [31:0] n1025;
  wire [3:0] n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire [3:0] n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire [33:0] n1036;
  wire xcsr_we;
  wire [11:0] xcsr_addr;
  wire [31:0] xcsr_wdata;
  wire [31:0] xcsr_rdata_pmp;
  wire [31:0] xcsr_rdata_alu;
  wire [31:0] xcsr_rdata_res;
  wire [31:0] xcsr_rdata_icc;
  wire clk_gated;
  wire [58:0] ctrl;
  wire [31:0] alu_imm;
  wire [31:0] rf_wdata;
  wire [31:0] rs1;
  wire [31:0] rs2;
  wire [31:0] rs3;
  wire [31:0] alu_res;
  wire [31:0] alu_add;
  wire [1:0] alu_cmp;
  wire [31:0] lsu_rdata;
  wire alu_cp_done;
  wire lsu_wait;
  wire [31:0] csr_rdata;
  wire [31:0] lsu_mar;
  wire [3:0] lsu_err;
  wire [31:0] pc_curr;
  wire [31:0] pc_ret;
  wire pmp_fault;
  wire [2:0] irq_machine;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[if_fence] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_wb_en] ;
  wire [4:0] \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rs1] ;
  wire [4:0] \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rs2] ;
  wire [4:0] \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rd] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_zero_we] ;
  wire [2:0] \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_op] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_sub] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_opa_mux] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_opb_mux] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_unsigned] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_alu] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_cfu] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_fpu] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_req] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_rw] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_mo_we] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_fence] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_priv] ;
  wire [2:0] \neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_funct3] ;
  wire [11:0] \neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_funct12] ;
  wire [6:0] \neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_opcode] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_priv] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_sleep] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_trap] ;
  wire \neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_debug] ;
  wire [31:0] \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[addr] ;
  wire [31:0] \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[data] ;
  wire [3:0] \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[ben] ;
  wire \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[stb] ;
  wire \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[rw] ;
  wire \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[src] ;
  wire \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[priv] ;
  wire \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[amo] ;
  wire [3:0] \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[amoop] ;
  wire \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[fence] ;
  wire \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[sleep] ;
  wire \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[debug] ;
  wire [31:0] \neorv32_cpu_control_inst.pc_next_o ;
  wire \neorv32_cpu_control_inst.xcsr_re_o ;
  wire [58:0] n1073;
  wire [79:0] n1075;
  wire [31:0] n1077;
  wire n1078;
  wire n1079;
  wire [1:0] n1089;
  wire [2:0] n1090;
  wire [31:0] n1091;
  wire [31:0] n1092;
  wire n1093;
  wire n1094;
  wire [4:0] n1095;
  wire [4:0] n1096;
  wire [4:0] n1097;
  wire n1098;
  wire [2:0] n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire [2:0] n1112;
  wire [11:0] n1113;
  wire [6:0] n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire [31:0] n1122;
  wire [31:0] n1123;
  wire [31:0] n1124;
  wire n1125;
  wire n1126;
  wire [4:0] n1127;
  wire [4:0] n1128;
  wire [4:0] n1129;
  wire n1130;
  wire [2:0] n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire [2:0] n1144;
  wire [11:0] n1145;
  wire [6:0] n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire [31:0] \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[addr] ;
  wire [31:0] \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[data] ;
  wire [3:0] \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[ben] ;
  wire \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[stb] ;
  wire \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[rw] ;
  wire \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[src] ;
  wire \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[priv] ;
  wire \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[amo] ;
  wire [3:0] \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[amoop] ;
  wire \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[fence] ;
  wire \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[sleep] ;
  wire \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[debug] ;
  wire n1156;
  wire n1157;
  wire [4:0] n1158;
  wire [4:0] n1159;
  wire [4:0] n1160;
  wire n1161;
  wire [2:0] n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire [2:0] n1175;
  wire [11:0] n1176;
  wire [6:0] n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire [79:0] n1186;
  wire [31:0] n1188;
  wire n1189;
  wire n1190;
  localparam [33:0] n1194 = 34'b0000000000000000000000000000000000;
  assign \icc_tx_o_icc_tx_o[rdy]  = n1005; //(module output)
  assign \icc_tx_o_icc_tx_o[ack]  = n1006; //(module output)
  assign \icc_tx_o_icc_tx_o[dat]  = n1007; //(module output)
  assign \ibus_req_o_ibus_req_o[addr]  = n1010; //(module output)
  assign \ibus_req_o_ibus_req_o[data]  = n1011; //(module output)
  assign \ibus_req_o_ibus_req_o[ben]  = n1012; //(module output)
  assign \ibus_req_o_ibus_req_o[stb]  = n1013; //(module output)
  assign \ibus_req_o_ibus_req_o[rw]  = n1014; //(module output)
  assign \ibus_req_o_ibus_req_o[src]  = n1015; //(module output)
  assign \ibus_req_o_ibus_req_o[priv]  = n1016; //(module output)
  assign \ibus_req_o_ibus_req_o[amo]  = n1017; //(module output)
  assign \ibus_req_o_ibus_req_o[amoop]  = n1018; //(module output)
  assign \ibus_req_o_ibus_req_o[fence]  = n1019; //(module output)
  assign \ibus_req_o_ibus_req_o[sleep]  = n1020; //(module output)
  assign \ibus_req_o_ibus_req_o[debug]  = n1021; //(module output)
  assign \dbus_req_o_dbus_req_o[addr]  = n1024; //(module output)
  assign \dbus_req_o_dbus_req_o[data]  = n1025; //(module output)
  assign \dbus_req_o_dbus_req_o[ben]  = n1026; //(module output)
  assign \dbus_req_o_dbus_req_o[stb]  = n1027; //(module output)
  assign \dbus_req_o_dbus_req_o[rw]  = n1028; //(module output)
  assign \dbus_req_o_dbus_req_o[src]  = n1029; //(module output)
  assign \dbus_req_o_dbus_req_o[priv]  = n1030; //(module output)
  assign \dbus_req_o_dbus_req_o[amo]  = n1031; //(module output)
  assign \dbus_req_o_dbus_req_o[amoop]  = n1032; //(module output)
  assign \dbus_req_o_dbus_req_o[fence]  = n1033; //(module output)
  assign \dbus_req_o_dbus_req_o[sleep]  = n1034; //(module output)
  assign \dbus_req_o_dbus_req_o[debug]  = n1035; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:712:12  */
  assign n1005 = n1194[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1026:14  */
  assign n1006 = n1194[1]; // extract
  assign n1007 = n1194[33:2]; // extract
  assign n1010 = n1075[31:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:711:12  */
  assign n1011 = n1075[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:122:3  */
  assign n1012 = n1075[67:64]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:124:5  */
  assign n1013 = n1075[68]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:124:5  */
  assign n1014 = n1075[69]; // extract
  assign n1015 = n1075[70]; // extract
  assign n1016 = n1075[71]; // extract
  assign n1017 = n1075[72]; // extract
  assign n1018 = n1075[76:73]; // extract
  assign n1019 = n1075[77]; // extract
  assign n1020 = n1075[78]; // extract
  assign n1021 = n1075[79]; // extract
  assign n1022 = {\ibus_rsp_i_ibus_rsp_i[err] , \ibus_rsp_i_ibus_rsp_i[ack] , \ibus_rsp_i_ibus_rsp_i[data] };
  assign n1024 = n1186[31:0]; // extract
  assign n1025 = n1186[63:32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:812:16  */
  assign n1026 = n1186[67:64]; // extract
  assign n1027 = n1186[68]; // extract
  assign n1028 = n1186[69]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:659:3  */
  assign n1029 = n1186[70]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:329:10  */
  assign n1030 = n1186[71]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:326:30  */
  assign n1031 = n1186[72]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:325:30  */
  assign n1032 = n1186[76:73]; // extract
  assign n1033 = n1186[77]; // extract
  assign n1034 = n1186[78]; // extract
  assign n1035 = n1186[79]; // extract
  assign n1036 = {\dbus_rsp_i_dbus_rsp_i[err] , \dbus_rsp_i_dbus_rsp_i[ack] , \dbus_rsp_i_dbus_rsp_i[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:109:10  */
  assign xcsr_rdata_pmp = 32'b00000000000000000000000000000000; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:111:10  */
  assign xcsr_rdata_res = n1092; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:112:10  */
  assign xcsr_rdata_icc = 32'b00000000000000000000000000000000; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:115:10  */
  assign clk_gated = clk_i; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:116:10  */
  assign ctrl = n1073; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:118:10  */
  assign rf_wdata = n1124; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:132:10  */
  assign pmp_fault = 1'b0; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:133:10  */
  assign irq_machine = n1090; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:213:3  */
  neorv32_cpu_control_0_1_40_d6061616ddd8e9e1dfd67ab5f4d47f4cb003c4e9 neorv32_cpu_control_inst (
    .clk_i(clk_gated),
    .clk_aux_i(clk_i),
    .rstn_i(rstn_i),
    .\ibus_rsp_i_ibus_rsp_i[data] (n1077),
    .\ibus_rsp_i_ibus_rsp_i[ack] (n1078),
    .\ibus_rsp_i_ibus_rsp_i[err] (n1079),
    .pmp_fault_i(pmp_fault),
    .alu_cp_done_i(alu_cp_done),
    .alu_cmp_i(alu_cmp),
    .alu_add_i(alu_add),
    .rf_rs1_i(rs1),
    .xcsr_rdata_i(xcsr_rdata_res),
    .irq_dbg_i(dbi_i),
    .irq_machine_i(irq_machine),
    .irq_fast_i(firq_i),
    .lsu_wait_i(lsu_wait),
    .lsu_mar_i(lsu_mar),
    .lsu_err_i(lsu_err),
    .\ctrl_o_ctrl_o[if_fence] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[if_fence] ),
    .\ctrl_o_ctrl_o[rf_wb_en] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_wb_en] ),
    .\ctrl_o_ctrl_o[rf_rs1] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rs1] ),
    .\ctrl_o_ctrl_o[rf_rs2] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rs2] ),
    .\ctrl_o_ctrl_o[rf_rd] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rd] ),
    .\ctrl_o_ctrl_o[rf_zero_we] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_zero_we] ),
    .\ctrl_o_ctrl_o[alu_op] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_op] ),
    .\ctrl_o_ctrl_o[alu_sub] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_sub] ),
    .\ctrl_o_ctrl_o[alu_opa_mux] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_opa_mux] ),
    .\ctrl_o_ctrl_o[alu_opb_mux] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_opb_mux] ),
    .\ctrl_o_ctrl_o[alu_unsigned] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_unsigned] ),
    .\ctrl_o_ctrl_o[alu_cp_alu] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_alu] ),
    .\ctrl_o_ctrl_o[alu_cp_cfu] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_cfu] ),
    .\ctrl_o_ctrl_o[alu_cp_fpu] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_fpu] ),
    .\ctrl_o_ctrl_o[lsu_req] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_req] ),
    .\ctrl_o_ctrl_o[lsu_rw] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_rw] ),
    .\ctrl_o_ctrl_o[lsu_mo_we] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_mo_we] ),
    .\ctrl_o_ctrl_o[lsu_fence] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_fence] ),
    .\ctrl_o_ctrl_o[lsu_priv] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_priv] ),
    .\ctrl_o_ctrl_o[ir_funct3] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_funct3] ),
    .\ctrl_o_ctrl_o[ir_funct12] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_funct12] ),
    .\ctrl_o_ctrl_o[ir_opcode] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_opcode] ),
    .\ctrl_o_ctrl_o[cpu_priv] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_priv] ),
    .\ctrl_o_ctrl_o[cpu_sleep] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_sleep] ),
    .\ctrl_o_ctrl_o[cpu_trap] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_trap] ),
    .\ctrl_o_ctrl_o[cpu_debug] (\neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_debug] ),
    .\ibus_req_o_ibus_req_o[addr] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[addr] ),
    .\ibus_req_o_ibus_req_o[data] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[data] ),
    .\ibus_req_o_ibus_req_o[ben] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[ben] ),
    .\ibus_req_o_ibus_req_o[stb] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[stb] ),
    .\ibus_req_o_ibus_req_o[rw] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[rw] ),
    .\ibus_req_o_ibus_req_o[src] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[src] ),
    .\ibus_req_o_ibus_req_o[priv] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[priv] ),
    .\ibus_req_o_ibus_req_o[amo] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[amo] ),
    .\ibus_req_o_ibus_req_o[amoop] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[amoop] ),
    .\ibus_req_o_ibus_req_o[fence] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[fence] ),
    .\ibus_req_o_ibus_req_o[sleep] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[sleep] ),
    .\ibus_req_o_ibus_req_o[debug] (\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[debug] ),
    .alu_imm_o(alu_imm),
    .pc_curr_o(pc_curr),
    .pc_next_o(),
    .pc_ret_o(pc_ret),
    .csr_rdata_o(csr_rdata),
    .xcsr_we_o(xcsr_we),
    .xcsr_re_o(),
    .xcsr_addr_o(xcsr_addr),
    .xcsr_wdata_o(xcsr_wdata));
  assign n1073 = {\neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_debug] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_trap] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_sleep] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[cpu_priv] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_opcode] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_funct12] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[ir_funct3] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_priv] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_fence] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_mo_we] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_rw] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[lsu_req] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_fpu] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_cfu] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_cp_alu] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_unsigned] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_opb_mux] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_opa_mux] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_sub] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[alu_op] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_zero_we] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rd] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rs2] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_rs1] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[rf_wb_en] , \neorv32_cpu_control_inst.ctrl_o_ctrl_o[if_fence] };
  assign n1075 = {\neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[debug] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[sleep] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[fence] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[amoop] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[amo] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[priv] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[src] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[rw] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[stb] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[ben] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[data] , \neorv32_cpu_control_inst.ibus_req_o_ibus_req_o[addr] };
  assign n1077 = n1022[31:0]; // extract
  assign n1078 = n1022[32]; // extract
  assign n1079 = n1022[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:298:24  */
  assign n1089 = {mti_i, mei_i};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:298:32  */
  assign n1090 = {n1089, msi_i};
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:301:36  */
  assign n1091 = xcsr_rdata_alu | xcsr_rdata_pmp;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:301:54  */
  assign n1092 = n1091 | xcsr_rdata_icc;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:306:3  */
  neorv32_cpu_regfile_9508e90548b0440a4a61e5743b76c1e309b23b7f neorv32_cpu_regfile_inst (
    .clk_i(clk_gated),
    .rstn_i(rstn_i),
    .\ctrl_i_ctrl_i[if_fence] (n1093),
    .\ctrl_i_ctrl_i[rf_wb_en] (n1094),
    .\ctrl_i_ctrl_i[rf_rs1] (n1095),
    .\ctrl_i_ctrl_i[rf_rs2] (n1096),
    .\ctrl_i_ctrl_i[rf_rd] (n1097),
    .\ctrl_i_ctrl_i[rf_zero_we] (n1098),
    .\ctrl_i_ctrl_i[alu_op] (n1099),
    .\ctrl_i_ctrl_i[alu_sub] (n1100),
    .\ctrl_i_ctrl_i[alu_opa_mux] (n1101),
    .\ctrl_i_ctrl_i[alu_opb_mux] (n1102),
    .\ctrl_i_ctrl_i[alu_unsigned] (n1103),
    .\ctrl_i_ctrl_i[alu_cp_alu] (n1104),
    .\ctrl_i_ctrl_i[alu_cp_cfu] (n1105),
    .\ctrl_i_ctrl_i[alu_cp_fpu] (n1106),
    .\ctrl_i_ctrl_i[lsu_req] (n1107),
    .\ctrl_i_ctrl_i[lsu_rw] (n1108),
    .\ctrl_i_ctrl_i[lsu_mo_we] (n1109),
    .\ctrl_i_ctrl_i[lsu_fence] (n1110),
    .\ctrl_i_ctrl_i[lsu_priv] (n1111),
    .\ctrl_i_ctrl_i[ir_funct3] (n1112),
    .\ctrl_i_ctrl_i[ir_funct12] (n1113),
    .\ctrl_i_ctrl_i[ir_opcode] (n1114),
    .\ctrl_i_ctrl_i[cpu_priv] (n1115),
    .\ctrl_i_ctrl_i[cpu_sleep] (n1116),
    .\ctrl_i_ctrl_i[cpu_trap] (n1117),
    .\ctrl_i_ctrl_i[cpu_debug] (n1118),
    .rd_i(rf_wdata),
    .rs1_o(rs1),
    .rs2_o(rs2),
    .rs3_o(rs3));
  assign n1093 = ctrl[0]; // extract
  assign n1094 = ctrl[1]; // extract
  assign n1095 = ctrl[6:2]; // extract
  assign n1096 = ctrl[11:7]; // extract
  assign n1097 = ctrl[16:12]; // extract
  assign n1098 = ctrl[17]; // extract
  assign n1099 = ctrl[20:18]; // extract
  assign n1100 = ctrl[21]; // extract
  assign n1101 = ctrl[22]; // extract
  assign n1102 = ctrl[23]; // extract
  assign n1103 = ctrl[24]; // extract
  assign n1104 = ctrl[25]; // extract
  assign n1105 = ctrl[26]; // extract
  assign n1106 = ctrl[27]; // extract
  assign n1107 = ctrl[28]; // extract
  assign n1108 = ctrl[29]; // extract
  assign n1109 = ctrl[30]; // extract
  assign n1110 = ctrl[31]; // extract
  assign n1111 = ctrl[32]; // extract
  assign n1112 = ctrl[35:33]; // extract
  assign n1113 = ctrl[47:36]; // extract
  assign n1114 = ctrl[54:48]; // extract
  assign n1115 = ctrl[55]; // extract
  assign n1116 = ctrl[56]; // extract
  assign n1117 = ctrl[57]; // extract
  assign n1118 = ctrl[58]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:325:23  */
  assign n1122 = alu_res | lsu_rdata;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:325:36  */
  assign n1123 = n1122 | csr_rdata;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:325:49  */
  assign n1124 = n1123 | pc_ret;
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:330:3  */
  neorv32_cpu_alu_f8bf199495d218f30da53ac11031539acc71c5ae neorv32_cpu_alu_inst (
    .clk_i(clk_gated),
    .rstn_i(rstn_i),
    .\ctrl_i_ctrl_i[if_fence] (n1125),
    .\ctrl_i_ctrl_i[rf_wb_en] (n1126),
    .\ctrl_i_ctrl_i[rf_rs1] (n1127),
    .\ctrl_i_ctrl_i[rf_rs2] (n1128),
    .\ctrl_i_ctrl_i[rf_rd] (n1129),
    .\ctrl_i_ctrl_i[rf_zero_we] (n1130),
    .\ctrl_i_ctrl_i[alu_op] (n1131),
    .\ctrl_i_ctrl_i[alu_sub] (n1132),
    .\ctrl_i_ctrl_i[alu_opa_mux] (n1133),
    .\ctrl_i_ctrl_i[alu_opb_mux] (n1134),
    .\ctrl_i_ctrl_i[alu_unsigned] (n1135),
    .\ctrl_i_ctrl_i[alu_cp_alu] (n1136),
    .\ctrl_i_ctrl_i[alu_cp_cfu] (n1137),
    .\ctrl_i_ctrl_i[alu_cp_fpu] (n1138),
    .\ctrl_i_ctrl_i[lsu_req] (n1139),
    .\ctrl_i_ctrl_i[lsu_rw] (n1140),
    .\ctrl_i_ctrl_i[lsu_mo_we] (n1141),
    .\ctrl_i_ctrl_i[lsu_fence] (n1142),
    .\ctrl_i_ctrl_i[lsu_priv] (n1143),
    .\ctrl_i_ctrl_i[ir_funct3] (n1144),
    .\ctrl_i_ctrl_i[ir_funct12] (n1145),
    .\ctrl_i_ctrl_i[ir_opcode] (n1146),
    .\ctrl_i_ctrl_i[cpu_priv] (n1147),
    .\ctrl_i_ctrl_i[cpu_sleep] (n1148),
    .\ctrl_i_ctrl_i[cpu_trap] (n1149),
    .\ctrl_i_ctrl_i[cpu_debug] (n1150),
    .csr_we_i(xcsr_we),
    .csr_addr_i(xcsr_addr),
    .csr_wdata_i(xcsr_wdata),
    .rs1_i(rs1),
    .rs2_i(rs2),
    .rs3_i(rs3),
    .pc_i(pc_curr),
    .imm_i(alu_imm),
    .csr_rdata_o(xcsr_rdata_alu),
    .cmp_o(alu_cmp),
    .res_o(alu_res),
    .add_o(alu_add),
    .cp_done_o(alu_cp_done));
  assign n1125 = ctrl[0]; // extract
  assign n1126 = ctrl[1]; // extract
  assign n1127 = ctrl[6:2]; // extract
  assign n1128 = ctrl[11:7]; // extract
  assign n1129 = ctrl[16:12]; // extract
  assign n1130 = ctrl[17]; // extract
  assign n1131 = ctrl[20:18]; // extract
  assign n1132 = ctrl[21]; // extract
  assign n1133 = ctrl[22]; // extract
  assign n1134 = ctrl[23]; // extract
  assign n1135 = ctrl[24]; // extract
  assign n1136 = ctrl[25]; // extract
  assign n1137 = ctrl[26]; // extract
  assign n1138 = ctrl[27]; // extract
  assign n1139 = ctrl[28]; // extract
  assign n1140 = ctrl[29]; // extract
  assign n1141 = ctrl[30]; // extract
  assign n1142 = ctrl[31]; // extract
  assign n1143 = ctrl[32]; // extract
  assign n1144 = ctrl[35:33]; // extract
  assign n1145 = ctrl[47:36]; // extract
  assign n1146 = ctrl[54:48]; // extract
  assign n1147 = ctrl[55]; // extract
  assign n1148 = ctrl[56]; // extract
  assign n1149 = ctrl[57]; // extract
  assign n1150 = ctrl[58]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_cpu.vhd:380:3  */
  neorv32_cpu_lsu_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_cpu_lsu_inst (
    .clk_i(clk_gated),
    .rstn_i(rstn_i),
    .\ctrl_i_ctrl_i[if_fence] (n1156),
    .\ctrl_i_ctrl_i[rf_wb_en] (n1157),
    .\ctrl_i_ctrl_i[rf_rs1] (n1158),
    .\ctrl_i_ctrl_i[rf_rs2] (n1159),
    .\ctrl_i_ctrl_i[rf_rd] (n1160),
    .\ctrl_i_ctrl_i[rf_zero_we] (n1161),
    .\ctrl_i_ctrl_i[alu_op] (n1162),
    .\ctrl_i_ctrl_i[alu_sub] (n1163),
    .\ctrl_i_ctrl_i[alu_opa_mux] (n1164),
    .\ctrl_i_ctrl_i[alu_opb_mux] (n1165),
    .\ctrl_i_ctrl_i[alu_unsigned] (n1166),
    .\ctrl_i_ctrl_i[alu_cp_alu] (n1167),
    .\ctrl_i_ctrl_i[alu_cp_cfu] (n1168),
    .\ctrl_i_ctrl_i[alu_cp_fpu] (n1169),
    .\ctrl_i_ctrl_i[lsu_req] (n1170),
    .\ctrl_i_ctrl_i[lsu_rw] (n1171),
    .\ctrl_i_ctrl_i[lsu_mo_we] (n1172),
    .\ctrl_i_ctrl_i[lsu_fence] (n1173),
    .\ctrl_i_ctrl_i[lsu_priv] (n1174),
    .\ctrl_i_ctrl_i[ir_funct3] (n1175),
    .\ctrl_i_ctrl_i[ir_funct12] (n1176),
    .\ctrl_i_ctrl_i[ir_opcode] (n1177),
    .\ctrl_i_ctrl_i[cpu_priv] (n1178),
    .\ctrl_i_ctrl_i[cpu_sleep] (n1179),
    .\ctrl_i_ctrl_i[cpu_trap] (n1180),
    .\ctrl_i_ctrl_i[cpu_debug] (n1181),
    .addr_i(alu_add),
    .wdata_i(rs2),
    .pmp_fault_i(pmp_fault),
    .\dbus_rsp_i_dbus_rsp_i[data] (n1188),
    .\dbus_rsp_i_dbus_rsp_i[ack] (n1189),
    .\dbus_rsp_i_dbus_rsp_i[err] (n1190),
    .rdata_o(lsu_rdata),
    .mar_o(lsu_mar),
    .wait_o(lsu_wait),
    .err_o(lsu_err),
    .\dbus_req_o_dbus_req_o[addr] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[addr] ),
    .\dbus_req_o_dbus_req_o[data] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[data] ),
    .\dbus_req_o_dbus_req_o[ben] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[ben] ),
    .\dbus_req_o_dbus_req_o[stb] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[stb] ),
    .\dbus_req_o_dbus_req_o[rw] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[rw] ),
    .\dbus_req_o_dbus_req_o[src] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[src] ),
    .\dbus_req_o_dbus_req_o[priv] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[priv] ),
    .\dbus_req_o_dbus_req_o[amo] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[amo] ),
    .\dbus_req_o_dbus_req_o[amoop] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[amoop] ),
    .\dbus_req_o_dbus_req_o[fence] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[fence] ),
    .\dbus_req_o_dbus_req_o[sleep] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[sleep] ),
    .\dbus_req_o_dbus_req_o[debug] (\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[debug] ));
  assign n1156 = ctrl[0]; // extract
  assign n1157 = ctrl[1]; // extract
  assign n1158 = ctrl[6:2]; // extract
  assign n1159 = ctrl[11:7]; // extract
  assign n1160 = ctrl[16:12]; // extract
  assign n1161 = ctrl[17]; // extract
  assign n1162 = ctrl[20:18]; // extract
  assign n1163 = ctrl[21]; // extract
  assign n1164 = ctrl[22]; // extract
  assign n1165 = ctrl[23]; // extract
  assign n1166 = ctrl[24]; // extract
  assign n1167 = ctrl[25]; // extract
  assign n1168 = ctrl[26]; // extract
  assign n1169 = ctrl[27]; // extract
  assign n1170 = ctrl[28]; // extract
  assign n1171 = ctrl[29]; // extract
  assign n1172 = ctrl[30]; // extract
  assign n1173 = ctrl[31]; // extract
  assign n1174 = ctrl[32]; // extract
  assign n1175 = ctrl[35:33]; // extract
  assign n1176 = ctrl[47:36]; // extract
  assign n1177 = ctrl[54:48]; // extract
  assign n1178 = ctrl[55]; // extract
  assign n1179 = ctrl[56]; // extract
  assign n1180 = ctrl[57]; // extract
  assign n1181 = ctrl[58]; // extract
  assign n1186 = {\neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[debug] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[sleep] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[fence] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[amoop] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[amo] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[priv] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[src] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[rw] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[stb] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[ben] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[data] , \neorv32_cpu_lsu_inst.dbus_req_o_dbus_req_o[addr] };
  assign n1188 = n1036[31:0]; // extract
  assign n1189 = n1036[32]; // extract
  assign n1190 = n1036[33]; // extract
endmodule

module neorv32_sys_clock_12
  (input  clk_i,
   input  rstn_i,
   input  [11:0] enable_i,
   output [7:0] clk_en_o);
  wire en;
  wire [11:0] cnt;
  wire [11:0] cnt2;
  wire n920;
  wire n928;
  wire n930;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire [11:0] n955;
  wire [11:0] n957;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  reg n1000;
  reg [11:0] n1001;
  reg [11:0] n1002;
  wire [7:0] n1003;
  assign clk_en_o = n1003; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:115:10  */
  assign en = n1000; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:116:10  */
  assign cnt = n1001; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:116:15  */
  assign cnt2 = n1002; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:124:16  */
  assign n920 = ~rstn_i;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n928 = enable_i[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n930 = 1'b0 | n928;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n932 = enable_i[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n933 = n930 | n932;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n934 = enable_i[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n935 = n933 | n934;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n936 = enable_i[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n937 = n935 | n936;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n938 = enable_i[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n939 = n937 | n938;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n940 = enable_i[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n941 = n939 | n940;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n942 = enable_i[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n943 = n941 | n942;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n944 = enable_i[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n945 = n943 | n944;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n946 = enable_i[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n947 = n945 | n946;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n948 = enable_i[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n949 = n947 | n948;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n950 = enable_i[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n951 = n949 | n950;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:30  */
  assign n952 = enable_i[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1030:22  */
  assign n953 = n951 | n952;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:131:48  */
  assign n955 = cnt + 12'b000000000001;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:130:7  */
  assign n957 = en ? n955 : 12'b000000000000;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:140:33  */
  assign n968 = cnt[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:140:51  */
  assign n969 = cnt2[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:140:43  */
  assign n970 = ~n969;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:140:38  */
  assign n971 = n968 & n970;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:141:33  */
  assign n972 = cnt[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:141:51  */
  assign n973 = cnt2[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:141:43  */
  assign n974 = ~n973;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:141:38  */
  assign n975 = n972 & n974;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:142:33  */
  assign n976 = cnt[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:142:51  */
  assign n977 = cnt2[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:142:43  */
  assign n978 = ~n977;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:142:38  */
  assign n979 = n976 & n978;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:143:33  */
  assign n980 = cnt[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:143:51  */
  assign n981 = cnt2[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:143:43  */
  assign n982 = ~n981;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:143:38  */
  assign n983 = n980 & n982;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:144:33  */
  assign n984 = cnt[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:144:51  */
  assign n985 = cnt2[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:144:43  */
  assign n986 = ~n985;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:144:38  */
  assign n987 = n984 & n986;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:145:33  */
  assign n988 = cnt[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:145:51  */
  assign n989 = cnt2[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:145:43  */
  assign n990 = ~n989;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:145:38  */
  assign n991 = n988 & n990;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:146:33  */
  assign n992 = cnt[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:146:51  */
  assign n993 = cnt2[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:146:43  */
  assign n994 = ~n993;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:146:38  */
  assign n995 = n992 & n994;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:147:33  */
  assign n996 = cnt[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:147:51  */
  assign n997 = cnt2[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:147:43  */
  assign n998 = ~n997;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:147:38  */
  assign n999 = n996 & n998;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:128:5  */
  always @(posedge clk_i or posedge n920)
    if (n920)
      n1000 <= 1'b0;
    else
      n1000 <= n953;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:128:5  */
  always @(posedge clk_i or posedge n920)
    if (n920)
      n1001 <= 12'b000000000000;
    else
      n1001 <= n957;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:128:5  */
  always @(posedge clk_i or posedge n920)
    if (n920)
      n1002 <= 12'b000000000000;
    else
      n1002 <= cnt;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:124:5  */
  assign n1003 = {n999, n995, n991, n987, n983, n979, n975, n971};
endmodule

module neorv32_sys_reset
  (input  clk_i,
   input  rstn_ext_i,
   input  rstn_wdt_i,
   input  rstn_dbg_i,
   output rstn_ext_o,
   output rstn_sys_o,
   output xrstn_wdt_o,
   output xrstn_ocd_o);
  wire [3:0] sreg_sys;
  wire [3:0] sreg_ext;
  wire n844;
  wire [2:0] n846;
  wire [3:0] n848;
  wire n855;
  wire n857;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire [2:0] n868;
  wire [3:0] n870;
  wire [3:0] n872;
  wire n879;
  wire n881;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n903;
  reg [3:0] n912;
  reg [3:0] n913;
  reg n914;
  reg n915;
  reg n916;
  reg n917;
  assign rstn_ext_o = n914; //(module output)
  assign rstn_sys_o = n915; //(module output)
  assign xrstn_wdt_o = n916; //(module output)
  assign xrstn_ocd_o = n917; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:36:10  */
  assign sreg_sys = n912; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:36:20  */
  assign sreg_ext = n913; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:44:20  */
  assign n844 = ~rstn_ext_i;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:51:29  */
  assign n846 = sreg_ext[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:51:56  */
  assign n848 = {n846, 1'b1};
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n855 = sreg_ext[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n857 = 1'b1 & n855;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n859 = sreg_ext[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n860 = n857 & n859;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n861 = sreg_ext[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n862 = n860 & n861;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n863 = sreg_ext[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n864 = n862 & n863;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:54:22  */
  assign n865 = ~rstn_wdt_i;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:54:44  */
  assign n866 = ~rstn_dbg_i;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:54:29  */
  assign n867 = n865 | n866;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:57:29  */
  assign n868 = sreg_sys[2:0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:57:56  */
  assign n870 = {n868, 1'b1};
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:54:7  */
  assign n872 = n867 ? 4'b0000 : n870;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n879 = sreg_sys[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n881 = 1'b1 & n879;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n883 = sreg_sys[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n884 = n881 & n883;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n885 = sreg_sys[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n886 = n884 & n885;
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:31  */
  assign n887 = sreg_sys[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_package.vhd:1042:22  */
  assign n888 = n886 & n887;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:68:20  */
  assign n903 = ~rstn_ext_i;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:49:5  */
  always @(posedge clk_i or posedge n844)
    if (n844)
      n912 <= 4'b0000;
    else
      n912 <= n872;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:49:5  */
  always @(posedge clk_i or posedge n844)
    if (n844)
      n913 <= 4'b0000;
    else
      n913 <= n848;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:49:5  */
  always @(posedge clk_i or posedge n844)
    if (n844)
      n914 <= 1'b0;
    else
      n914 <= n864;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:49:5  */
  always @(posedge clk_i or posedge n844)
    if (n844)
      n915 <= 1'b0;
    else
      n915 <= n888;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:71:5  */
  always @(posedge clk_i or posedge n903)
    if (n903)
      n916 <= 1'b0;
    else
      n916 <= rstn_wdt_i;
  /* ../../ext/neorv32/rtl/core/neorv32_sys.vhd:71:5  */
  always @(posedge clk_i or posedge n903)
    if (n903)
      n917 <= 1'b0;
    else
      n917 <= rstn_dbg_i;
endmodule

module neorv32_top_98304000_0_0_4_1_40_16384_16384_4_64_4_64_255_64_32_16_64_23_1_1_1_1_1_1_1_1_2_1_32_32_1_1_1_1_14ddc86578158058671fcea0fd4647c83d242e3e
  (input  clk_i,
   input  rstn_i,
   input  jtag_tck_i,
   input  jtag_tdi_i,
   input  jtag_tms_i,
   input  jtagspi_sdi_i,
   input  [31:0] xbus_dat_i,
   input  xbus_ack_i,
   input  xbus_err_i,
   input  [31:0] slink_rx_dat_i,
   input  [3:0] slink_rx_src_i,
   input  slink_rx_val_i,
   input  slink_rx_lst_i,
   input  slink_tx_rdy_i,
   input  xip_dat_i,
   input  [31:0] gpio_i,
   input  uart0_rxd_i,
   input  uart0_cts_i,
   input  uart1_rxd_i,
   input  uart1_cts_i,
   input  spi_dat_i,
   input  sdi_clk_i,
   input  sdi_dat_i,
   input  sdi_csn_i,
   input  twi_sda_i,
   input  twi_scl_i,
   input  twd_sda_i,
   input  twd_scl_i,
   input  onewire_i,
   input  [31:0] cfs_in_i,
   input  mtime_irq_i,
   input  msw_irq_i,
   input  mext_irq_i,
   output rstn_ocd_o,
   output rstn_wdt_o,
   output jtag_tdo_o,
   output jtagspi_sck_o,
   output jtagspi_sdo_o,
   output jtagspi_csn_o,
   output [31:0] xbus_adr_o,
   output [31:0] xbus_dat_o,
   output [2:0] xbus_tag_o,
   output xbus_we_o,
   output [3:0] xbus_sel_o,
   output xbus_stb_o,
   output xbus_cyc_o,
   output slink_rx_rdy_o,
   output [31:0] slink_tx_dat_o,
   output [3:0] slink_tx_dst_o,
   output slink_tx_val_o,
   output slink_tx_lst_o,
   output xip_csn_o,
   output xip_clk_o,
   output xip_dat_o,
   output [31:0] gpio_o,
   output uart0_txd_o,
   output uart0_rts_o,
   output uart1_txd_o,
   output uart1_rts_o,
   output spi_clk_o,
   output spi_dat_o,
   output [7:0] spi_csn_o,
   output sdi_dat_o,
   output twi_sda_o,
   output twi_scl_o,
   output twd_sda_o,
   output twd_scl_o,
   output onewire_o,
   output [15:0] pwm_o,
   output [31:0] cfs_out_o,
   output neoled_o,
   output [63:0] mtime_time_o);
  wire rstn_wdt;
  wire rstn_sys;
  wire rstn_ext;
  wire [7:0] clk_gen;
  wire [11:0] clk_gen_en;
  wire [11:0] clk_gen_en2;
  wire [40:0] dmi_req;
  wire [32:0] dmi_rsp;
  wire dci_ndmrstn;
  wire dci_haltreq;
  wire [33:0] icc_tx;
  wire [33:0] icc_rx;
  wire [79:0] cpu_i_req;
  wire [79:0] cpu_d_req;
  wire [79:0] icache_req;
  wire [79:0] dcache_req;
  wire [79:0] core_req;
  wire [33:0] cpu_i_rsp;
  wire [33:0] cpu_d_rsp;
  wire [33:0] icache_rsp;
  wire [33:0] dcache_rsp;
  wire [33:0] core_rsp;
  wire [79:0] sys1_req;
  wire [79:0] sys2_req;
  wire [79:0] sys3_req;
  wire [33:0] sys1_rsp;
  wire [33:0] sys2_rsp;
  wire [33:0] sys3_rsp;
  wire [79:0] dmem_req;
  wire [79:0] xipcache_req;
  wire [79:0] xip_req;
  wire [79:0] io_req;
  wire [79:0] xcache_req;
  wire [79:0] xbus_req;
  wire [33:0] imem_rsp;
  wire [33:0] dmem_rsp;
  wire [33:0] xipcache_rsp;
  wire [33:0] xip_rsp;
  wire [33:0] io_rsp;
  wire [33:0] xcache_rsp;
  wire [33:0] xbus_rsp;
  wire [1759:0] iodev_req;
  wire [747:0] iodev_rsp;
  wire [15:0] firq;
  wire [15:0] cpu_firq;
  wire mtime_irq;
  wire msw_irq;
  wire \soc_generators_neorv32_sys_reset_inst.xrstn_wdt_o ;
  wire \soc_generators_neorv32_sys_reset_inst.xrstn_ocd_o ;
  wire n225;
  wire n226;
  wire [1:0] n227;
  wire n228;
  wire [2:0] n229;
  wire n230;
  wire [3:0] n231;
  wire n232;
  wire [4:0] n233;
  wire n234;
  wire [5:0] n235;
  wire n236;
  wire [6:0] n237;
  wire n238;
  wire [7:0] n239;
  wire n240;
  wire [8:0] n241;
  wire n242;
  wire [9:0] n243;
  wire n244;
  wire [10:0] n245;
  wire n246;
  wire [11:0] n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire \core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[rdy] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[ack] ;
  wire [31:0] \core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[dat] ;
  wire [31:0] \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[addr] ;
  wire [31:0] \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[data] ;
  wire [3:0] \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[ben] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[stb] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[rw] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[src] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[priv] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[amo] ;
  wire [3:0] \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[amoop] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[fence] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[sleep] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[debug] ;
  wire [31:0] \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[addr] ;
  wire [31:0] \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[data] ;
  wire [3:0] \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[ben] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[stb] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[rw] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[src] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[priv] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[amo] ;
  wire [3:0] \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[amoop] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[fence] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[sleep] ;
  wire \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[debug] ;
  wire [33:0] n264;
  wire n266;
  wire n267;
  wire [31:0] n268;
  wire [79:0] n269;
  wire [31:0] n271;
  wire n272;
  wire n273;
  wire [79:0] n274;
  wire [31:0] n276;
  wire n277;
  wire n278;
  wire [31:0] \core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[data] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[ack] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[err] ;
  wire [31:0] \core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[data] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[ack] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[err] ;
  wire [31:0] \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[addr] ;
  wire [31:0] \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[data] ;
  wire [3:0] \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[ben] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[stb] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[rw] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[src] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[priv] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[amo] ;
  wire [3:0] \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[amoop] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[fence] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[sleep] ;
  wire \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[debug] ;
  localparam n279 = 1'b0;
  wire [31:0] n280;
  wire [31:0] n281;
  wire [3:0] n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire [3:0] n288;
  wire n289;
  wire n290;
  wire n291;
  wire [33:0] n292;
  wire [31:0] n294;
  wire [31:0] n295;
  wire [3:0] n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire [3:0] n302;
  wire n303;
  wire n304;
  wire n305;
  wire [33:0] n306;
  wire [79:0] n308;
  wire [31:0] n310;
  wire n311;
  wire n312;
  localparam [33:0] n315 = 34'b0000000000000000000000000000000000;
  wire [31:0] \neorv32_bus_gateway_inst.rsp_o_rsp_o[data] ;
  wire \neorv32_bus_gateway_inst.rsp_o_rsp_o[ack] ;
  wire \neorv32_bus_gateway_inst.rsp_o_rsp_o[err] ;
  wire [31:0] \neorv32_bus_gateway_inst.a_req_o_a_req_o[addr] ;
  wire [31:0] \neorv32_bus_gateway_inst.a_req_o_a_req_o[data] ;
  wire [3:0] \neorv32_bus_gateway_inst.a_req_o_a_req_o[ben] ;
  wire \neorv32_bus_gateway_inst.a_req_o_a_req_o[stb] ;
  wire \neorv32_bus_gateway_inst.a_req_o_a_req_o[rw] ;
  wire \neorv32_bus_gateway_inst.a_req_o_a_req_o[src] ;
  wire \neorv32_bus_gateway_inst.a_req_o_a_req_o[priv] ;
  wire \neorv32_bus_gateway_inst.a_req_o_a_req_o[amo] ;
  wire [3:0] \neorv32_bus_gateway_inst.a_req_o_a_req_o[amoop] ;
  wire \neorv32_bus_gateway_inst.a_req_o_a_req_o[fence] ;
  wire \neorv32_bus_gateway_inst.a_req_o_a_req_o[sleep] ;
  wire \neorv32_bus_gateway_inst.a_req_o_a_req_o[debug] ;
  wire [31:0] \neorv32_bus_gateway_inst.b_req_o_b_req_o[addr] ;
  wire [31:0] \neorv32_bus_gateway_inst.b_req_o_b_req_o[data] ;
  wire [3:0] \neorv32_bus_gateway_inst.b_req_o_b_req_o[ben] ;
  wire \neorv32_bus_gateway_inst.b_req_o_b_req_o[stb] ;
  wire \neorv32_bus_gateway_inst.b_req_o_b_req_o[rw] ;
  wire \neorv32_bus_gateway_inst.b_req_o_b_req_o[src] ;
  wire \neorv32_bus_gateway_inst.b_req_o_b_req_o[priv] ;
  wire \neorv32_bus_gateway_inst.b_req_o_b_req_o[amo] ;
  wire [3:0] \neorv32_bus_gateway_inst.b_req_o_b_req_o[amoop] ;
  wire \neorv32_bus_gateway_inst.b_req_o_b_req_o[fence] ;
  wire \neorv32_bus_gateway_inst.b_req_o_b_req_o[sleep] ;
  wire \neorv32_bus_gateway_inst.b_req_o_b_req_o[debug] ;
  wire [31:0] \neorv32_bus_gateway_inst.c_req_o_c_req_o[addr] ;
  wire [31:0] \neorv32_bus_gateway_inst.c_req_o_c_req_o[data] ;
  wire [3:0] \neorv32_bus_gateway_inst.c_req_o_c_req_o[ben] ;
  wire \neorv32_bus_gateway_inst.c_req_o_c_req_o[stb] ;
  wire \neorv32_bus_gateway_inst.c_req_o_c_req_o[rw] ;
  wire \neorv32_bus_gateway_inst.c_req_o_c_req_o[src] ;
  wire \neorv32_bus_gateway_inst.c_req_o_c_req_o[priv] ;
  wire \neorv32_bus_gateway_inst.c_req_o_c_req_o[amo] ;
  wire [3:0] \neorv32_bus_gateway_inst.c_req_o_c_req_o[amoop] ;
  wire \neorv32_bus_gateway_inst.c_req_o_c_req_o[fence] ;
  wire \neorv32_bus_gateway_inst.c_req_o_c_req_o[sleep] ;
  wire \neorv32_bus_gateway_inst.c_req_o_c_req_o[debug] ;
  wire [31:0] \neorv32_bus_gateway_inst.d_req_o_d_req_o[addr] ;
  wire [31:0] \neorv32_bus_gateway_inst.d_req_o_d_req_o[data] ;
  wire [3:0] \neorv32_bus_gateway_inst.d_req_o_d_req_o[ben] ;
  wire \neorv32_bus_gateway_inst.d_req_o_d_req_o[stb] ;
  wire \neorv32_bus_gateway_inst.d_req_o_d_req_o[rw] ;
  wire \neorv32_bus_gateway_inst.d_req_o_d_req_o[src] ;
  wire \neorv32_bus_gateway_inst.d_req_o_d_req_o[priv] ;
  wire \neorv32_bus_gateway_inst.d_req_o_d_req_o[amo] ;
  wire [3:0] \neorv32_bus_gateway_inst.d_req_o_d_req_o[amoop] ;
  wire \neorv32_bus_gateway_inst.d_req_o_d_req_o[fence] ;
  wire \neorv32_bus_gateway_inst.d_req_o_d_req_o[sleep] ;
  wire \neorv32_bus_gateway_inst.d_req_o_d_req_o[debug] ;
  wire [31:0] \neorv32_bus_gateway_inst.x_req_o_x_req_o[addr] ;
  wire [31:0] \neorv32_bus_gateway_inst.x_req_o_x_req_o[data] ;
  wire [3:0] \neorv32_bus_gateway_inst.x_req_o_x_req_o[ben] ;
  wire \neorv32_bus_gateway_inst.x_req_o_x_req_o[stb] ;
  wire \neorv32_bus_gateway_inst.x_req_o_x_req_o[rw] ;
  wire \neorv32_bus_gateway_inst.x_req_o_x_req_o[src] ;
  wire \neorv32_bus_gateway_inst.x_req_o_x_req_o[priv] ;
  wire \neorv32_bus_gateway_inst.x_req_o_x_req_o[amo] ;
  wire [3:0] \neorv32_bus_gateway_inst.x_req_o_x_req_o[amoop] ;
  wire \neorv32_bus_gateway_inst.x_req_o_x_req_o[fence] ;
  wire \neorv32_bus_gateway_inst.x_req_o_x_req_o[sleep] ;
  wire \neorv32_bus_gateway_inst.x_req_o_x_req_o[debug] ;
  wire [31:0] n317;
  wire [31:0] n318;
  wire [3:0] n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire [3:0] n325;
  wire n326;
  wire n327;
  wire n328;
  wire [33:0] n329;
  wire [31:0] n333;
  wire n334;
  wire n335;
  wire [79:0] n336;
  wire [31:0] n338;
  wire n339;
  wire n340;
  wire [79:0] n341;
  wire [31:0] n343;
  wire n344;
  wire n345;
  wire [79:0] n346;
  wire [31:0] n348;
  wire n349;
  wire n350;
  wire [79:0] n351;
  wire [31:0] n353;
  wire n354;
  wire n355;
  wire [31:0] \memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire [31:0] n357;
  wire [31:0] n358;
  wire [3:0] n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire [3:0] n365;
  wire n366;
  wire n367;
  wire n368;
  wire [33:0] n369;
  wire [31:0] \memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire [31:0] \memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[data] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[ack] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[err] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xip_inst.clkgen_en_o ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_csn_o ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_clk_o ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_dat_o ;
  wire [79:0] n371;
  wire [31:0] n372;
  wire [31:0] n373;
  wire [3:0] n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire [3:0] n380;
  wire n381;
  wire n382;
  wire n383;
  wire [33:0] n384;
  wire [31:0] n386;
  wire [31:0] n387;
  wire [3:0] n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire [3:0] n394;
  wire n395;
  wire n396;
  wire n397;
  wire [33:0] n398;
  wire [31:0] \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[data] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[ack] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[err] ;
  wire [31:0] \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[addr] ;
  wire [31:0] \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[data] ;
  wire [3:0] \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[ben] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[stb] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[rw] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[src] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[priv] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[amo] ;
  wire [3:0] \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[amoop] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[fence] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[sleep] ;
  wire \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[debug] ;
  wire [31:0] n404;
  wire [31:0] n405;
  wire [3:0] n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire [3:0] n412;
  wire n413;
  wire n414;
  wire n415;
  wire [33:0] n416;
  wire [79:0] n418;
  wire [31:0] n420;
  wire n421;
  wire n422;
  wire [31:0] \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire [31:0] \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_adr_o ;
  wire [31:0] \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_dat_o ;
  wire [2:0] \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_tag_o ;
  wire \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_we_o ;
  wire [3:0] \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_sel_o ;
  wire \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_stb_o ;
  wire \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_cyc_o ;
  wire [31:0] n423;
  wire [31:0] n424;
  wire [3:0] n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire [3:0] n431;
  wire n432;
  wire n433;
  wire n434;
  wire [33:0] n435;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[data] ;
  wire \io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[ack] ;
  wire \io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[err] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_01_req_o_dev_01_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_02_req_o_dev_02_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_03_req_o_dev_03_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_04_req_o_dev_04_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_05_req_o_dev_05_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_06_req_o_dev_06_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_07_req_o_dev_07_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_08_req_o_dev_08_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_09_req_o_dev_09_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_19_req_o_dev_19_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[debug] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[addr] ;
  wire [31:0] \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[data] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[ben] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[stb] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[rw] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[src] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[priv] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[amo] ;
  wire [3:0] \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[amoop] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[fence] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[sleep] ;
  wire \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[debug] ;
  wire [31:0] n444;
  wire [31:0] n445;
  wire [3:0] n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire [3:0] n452;
  wire n453;
  wire n454;
  wire n455;
  wire [33:0] n456;
  wire [79:0] n458;
  wire [33:0] n460;
  wire [31:0] n461;
  wire n462;
  wire n463;
  wire [31:0] n465;
  wire n466;
  wire n467;
  wire [31:0] n469;
  wire n470;
  wire n471;
  wire [31:0] n473;
  wire n474;
  wire n475;
  wire [31:0] n477;
  wire n478;
  wire n479;
  wire [31:0] n481;
  wire n482;
  wire n483;
  wire [31:0] n485;
  wire n486;
  wire n487;
  wire [31:0] n489;
  wire n490;
  wire n491;
  wire [31:0] n493;
  wire n494;
  wire n495;
  wire [31:0] n497;
  wire n498;
  wire n499;
  wire [79:0] n500;
  wire [33:0] n502;
  wire [31:0] n503;
  wire n504;
  wire n505;
  wire [79:0] n506;
  wire [33:0] n508;
  wire [31:0] n509;
  wire n510;
  wire n511;
  wire [79:0] n512;
  wire [33:0] n514;
  wire [31:0] n515;
  wire n516;
  wire n517;
  wire [79:0] n518;
  wire [33:0] n520;
  wire [31:0] n521;
  wire n522;
  wire n523;
  wire [79:0] n524;
  wire [33:0] n526;
  wire [31:0] n527;
  wire n528;
  wire n529;
  wire [79:0] n530;
  wire [33:0] n532;
  wire [31:0] n533;
  wire n534;
  wire n535;
  wire [79:0] n536;
  wire [33:0] n538;
  wire [31:0] n539;
  wire n540;
  wire n541;
  wire [79:0] n542;
  wire [33:0] n544;
  wire [31:0] n545;
  wire n546;
  wire n547;
  wire [79:0] n548;
  wire [33:0] n550;
  wire [31:0] n551;
  wire n552;
  wire n553;
  wire [31:0] n555;
  wire n556;
  wire n557;
  wire [79:0] n558;
  wire [33:0] n560;
  wire [31:0] n561;
  wire n562;
  wire n563;
  wire [79:0] n564;
  wire [33:0] n566;
  wire [31:0] n567;
  wire n568;
  wire n569;
  wire [79:0] n570;
  wire [33:0] n572;
  wire [31:0] n573;
  wire n574;
  wire n575;
  wire [79:0] n576;
  wire [33:0] n578;
  wire [31:0] n579;
  wire n580;
  wire n581;
  wire [79:0] n582;
  wire [33:0] n584;
  wire [31:0] n585;
  wire n586;
  wire n587;
  wire [79:0] n588;
  wire [33:0] n590;
  wire [31:0] n591;
  wire n592;
  wire n593;
  wire [79:0] n594;
  wire [33:0] n596;
  wire [31:0] n597;
  wire n598;
  wire n599;
  wire [79:0] n600;
  wire [33:0] n602;
  wire [31:0] n603;
  wire n604;
  wire n605;
  wire [79:0] n606;
  wire [33:0] n608;
  wire [31:0] n609;
  wire n610;
  wire n611;
  wire [79:0] n612;
  wire [33:0] n614;
  wire [31:0] n615;
  wire n616;
  wire n617;
  wire [79:0] n618;
  wire [33:0] n620;
  wire [31:0] n621;
  wire n622;
  wire n623;
  wire [79:0] n624;
  wire [33:0] n626;
  wire [31:0] n627;
  wire n628;
  wire n629;
  wire [31:0] \io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire [79:0] n630;
  wire [31:0] n631;
  wire [31:0] n632;
  wire [3:0] n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire [3:0] n639;
  wire n640;
  wire n641;
  wire n642;
  wire [33:0] n643;
  localparam [31:0] n647 = 32'b00000000000000000000000000000000;
  localparam n648 = 1'b0;
  wire [31:0] \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire [31:0] \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.gpio_o ;
  wire \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.cpu_irq_o ;
  wire [79:0] n650;
  wire [31:0] n651;
  wire [31:0] n652;
  wire [3:0] n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire [3:0] n659;
  wire n660;
  wire n661;
  wire n662;
  wire [33:0] n663;
  wire [31:0] \io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire [63:0] \io_system_neorv32_clint_enabled_neorv32_clint_inst.time_o ;
  wire [79:0] n669;
  wire [31:0] n670;
  wire [31:0] n671;
  wire [3:0] n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire [3:0] n678;
  wire n679;
  wire n680;
  wire n681;
  wire [33:0] n682;
  wire [31:0] \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.clkgen_en_o ;
  wire \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.uart_txd_o ;
  wire \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.uart_rts_o ;
  wire \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.irq_rx_o ;
  wire \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.irq_tx_o ;
  wire [79:0] n687;
  wire [31:0] n688;
  wire [31:0] n689;
  wire [3:0] n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire [3:0] n696;
  wire n697;
  wire n698;
  wire n699;
  wire [33:0] n700;
  localparam n707 = 1'b0;
  localparam n708 = 1'b1;
  wire [31:0] \io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire \io_system_neorv32_spi_enabled_neorv32_spi_inst.clkgen_en_o ;
  wire \io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_clk_o ;
  wire \io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_dat_o ;
  wire [7:0] \io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_csn_o ;
  wire \io_system_neorv32_spi_enabled_neorv32_spi_inst.irq_o ;
  wire [79:0] n712;
  wire [31:0] n713;
  wire [31:0] n714;
  wire [3:0] n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire [3:0] n721;
  wire n722;
  wire n723;
  wire n724;
  wire [33:0] n725;
  wire [31:0] \io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire \io_system_neorv32_twi_enabled_neorv32_twi_inst.clkgen_en_o ;
  wire \io_system_neorv32_twi_enabled_neorv32_twi_inst.twi_sda_o ;
  wire \io_system_neorv32_twi_enabled_neorv32_twi_inst.twi_scl_o ;
  wire \io_system_neorv32_twi_enabled_neorv32_twi_inst.irq_o ;
  wire [79:0] n732;
  wire [31:0] n733;
  wire [31:0] n734;
  wire [3:0] n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire [3:0] n741;
  wire n742;
  wire n743;
  wire n744;
  wire [33:0] n745;
  localparam n751 = 1'b1;
  localparam n752 = 1'b1;
  wire [31:0] \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.clkgen_en_o ;
  wire [15:0] \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.pwm_o ;
  wire [79:0] n755;
  wire [31:0] n756;
  wire [31:0] n757;
  wire [3:0] n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire [3:0] n764;
  wire n765;
  wire n766;
  wire n767;
  wire [33:0] n768;
  localparam n774 = 1'b0;
  localparam n777 = 1'b1;
  localparam n782 = 1'b0;
  localparam [31:0] n783 = 32'b00000000000000000000000000000000;
  localparam [3:0] n784 = 4'b0000;
  localparam n785 = 1'b0;
  localparam n786 = 1'b0;
  wire [31:0] \io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire [79:0] n787;
  wire [31:0] n788;
  wire [31:0] n789;
  wire [3:0] n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire [3:0] n796;
  wire n797;
  wire n798;
  wire n799;
  wire [33:0] n800;
  wire \neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtag_tdo_o ;
  wire [6:0] \neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[addr] ;
  wire [1:0] \neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[op] ;
  wire [31:0] \neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[data] ;
  wire \neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_sck_o ;
  wire \neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_sdo_o ;
  wire \neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_csn_o ;
  wire [40:0] n803;
  wire [31:0] n805;
  wire n806;
  wire [31:0] \neorv32_ocd_enabled_neorv32_debug_dm_inst.dmi_rsp_o_dmi_rsp_o[data] ;
  wire \neorv32_ocd_enabled_neorv32_debug_dm_inst.dmi_rsp_o_dmi_rsp_o[ack] ;
  wire [31:0] \neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[data] ;
  wire \neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[ack] ;
  wire \neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[err] ;
  wire [6:0] n810;
  wire [1:0] n811;
  wire [31:0] n812;
  wire [32:0] n813;
  wire [79:0] n815;
  wire [31:0] n816;
  wire [31:0] n817;
  wire [3:0] n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire [3:0] n824;
  wire n825;
  wire n826;
  wire n827;
  wire [33:0] n828;
  wire [11:0] n832;
  wire [1759:0] n835;
  wire [747:0] n836;
  wire [15:0] n837;
  wire [15:0] n838;
  assign rstn_ocd_o = \soc_generators_neorv32_sys_reset_inst.xrstn_ocd_o ; //(module output)
  assign rstn_wdt_o = \soc_generators_neorv32_sys_reset_inst.xrstn_wdt_o ; //(module output)
  assign jtag_tdo_o = \neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtag_tdo_o ; //(module output)
  assign jtagspi_sck_o = \neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_sck_o ; //(module output)
  assign jtagspi_sdo_o = \neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_sdo_o ; //(module output)
  assign jtagspi_csn_o = \neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_csn_o ; //(module output)
  assign xbus_adr_o = \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_adr_o ; //(module output)
  assign xbus_dat_o = \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_dat_o ; //(module output)
  assign xbus_tag_o = \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_tag_o ; //(module output)
  assign xbus_we_o = \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_we_o ; //(module output)
  assign xbus_sel_o = \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_sel_o ; //(module output)
  assign xbus_stb_o = \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_stb_o ; //(module output)
  assign xbus_cyc_o = \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_cyc_o ; //(module output)
  assign slink_rx_rdy_o = n782; //(module output)
  assign slink_tx_dat_o = n783; //(module output)
  assign slink_tx_dst_o = n784; //(module output)
  assign slink_tx_val_o = n785; //(module output)
  assign slink_tx_lst_o = n786; //(module output)
  assign xip_csn_o = \memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_csn_o ; //(module output)
  assign xip_clk_o = \memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_clk_o ; //(module output)
  assign xip_dat_o = \memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_dat_o ; //(module output)
  assign gpio_o = \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.gpio_o ; //(module output)
  assign uart0_txd_o = \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.uart_txd_o ; //(module output)
  assign uart0_rts_o = \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.uart_rts_o ; //(module output)
  assign uart1_txd_o = n707; //(module output)
  assign uart1_rts_o = n708; //(module output)
  assign spi_clk_o = \io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_clk_o ; //(module output)
  assign spi_dat_o = \io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_dat_o ; //(module output)
  assign spi_csn_o = \io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_csn_o ; //(module output)
  assign sdi_dat_o = n648; //(module output)
  assign twi_sda_o = \io_system_neorv32_twi_enabled_neorv32_twi_inst.twi_sda_o ; //(module output)
  assign twi_scl_o = \io_system_neorv32_twi_enabled_neorv32_twi_inst.twi_scl_o ; //(module output)
  assign twd_sda_o = n751; //(module output)
  assign twd_scl_o = n752; //(module output)
  assign onewire_o = n777; //(module output)
  assign pwm_o = \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.pwm_o ; //(module output)
  assign cfs_out_o = n647; //(module output)
  assign neoled_o = n774; //(module output)
  assign mtime_time_o = \io_system_neorv32_clint_enabled_neorv32_clint_inst.time_o ; //(module output)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:294:10  */
  assign rstn_wdt = 1'b1; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:303:10  */
  assign clk_gen_en = n832; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:304:10  */
  assign clk_gen_en2 = n247; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:307:10  */
  assign dmi_req = n803; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:308:10  */
  assign dmi_rsp = n813; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:316:10  */
  assign icc_tx = n264; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:316:18  */
  assign icc_rx = icc_tx; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:321:10  */
  assign cpu_i_req = n269; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:321:21  */
  assign cpu_d_req = n274; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:321:32  */
  assign icache_req = cpu_i_req; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:321:44  */
  assign dcache_req = cpu_d_req; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:321:56  */
  assign core_req = n308; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:322:10  */
  assign cpu_i_rsp = icache_rsp; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:322:21  */
  assign cpu_d_rsp = dcache_rsp; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:322:32  */
  assign icache_rsp = n306; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:322:44  */
  assign dcache_rsp = n292; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:322:56  */
  assign core_rsp = sys1_rsp; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:325:10  */
  assign sys1_req = core_req; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:325:20  */
  assign sys2_req = sys1_req; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:325:39  */
  assign sys3_req = sys2_req; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:326:10  */
  assign sys1_rsp = sys2_rsp; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:326:20  */
  assign sys2_rsp = sys3_rsp; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:326:39  */
  assign sys3_rsp = n329; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:329:20  */
  assign dmem_req = n336; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:329:30  */
  assign xipcache_req = n418; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:329:44  */
  assign xip_req = n341; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:329:53  */
  assign io_req = n346; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:329:61  */
  assign xcache_req = xbus_req; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:329:73  */
  assign xbus_req = n351; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:330:10  */
  assign imem_rsp = 34'b0000000000000000000000000000000000; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:330:20  */
  assign dmem_rsp = n369; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:330:30  */
  assign xipcache_rsp = n398; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:330:44  */
  assign xip_rsp = n416; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:330:53  */
  assign io_rsp = n456; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:330:61  */
  assign xcache_rsp = n435; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:330:73  */
  assign xbus_rsp = xcache_rsp; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:340:10  */
  assign iodev_req = n835; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:341:10  */
  assign iodev_rsp = n836; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:349:10  */
  assign firq = n837; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:350:10  */
  assign cpu_firq = n838; // (signal)
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:443:5  */
  neorv32_sys_reset soc_generators_neorv32_sys_reset_inst (
    .clk_i(clk_i),
    .rstn_ext_i(rstn_i),
    .rstn_wdt_i(rstn_wdt),
    .rstn_dbg_i(dci_ndmrstn),
    .rstn_ext_o(rstn_ext),
    .rstn_sys_o(rstn_sys),
    .xrstn_wdt_o(\soc_generators_neorv32_sys_reset_inst.xrstn_wdt_o ),
    .xrstn_ocd_o(\soc_generators_neorv32_sys_reset_inst.xrstn_ocd_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:458:5  */
  neorv32_sys_clock_12 soc_generators_neorv32_sys_clock_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .enable_i(clk_gen_en2),
    .clk_en_o(clk_gen));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:470:30  */
  assign n225 = clk_gen_en[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:470:54  */
  assign n226 = clk_gen_en[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:470:42  */
  assign n227 = {n225, n226};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:470:77  */
  assign n228 = clk_gen_en[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:470:65  */
  assign n229 = {n227, n228};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:470:100  */
  assign n230 = clk_gen_en[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:470:88  */
  assign n231 = {n229, n230};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:471:30  */
  assign n232 = clk_gen_en[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:470:109  */
  assign n233 = {n231, n232};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:471:54  */
  assign n234 = clk_gen_en[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:471:42  */
  assign n235 = {n233, n234};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:471:77  */
  assign n236 = clk_gen_en[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:471:65  */
  assign n237 = {n235, n236};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:471:100  */
  assign n238 = clk_gen_en[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:471:88  */
  assign n239 = {n237, n238};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:472:30  */
  assign n240 = clk_gen_en[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:471:109  */
  assign n241 = {n239, n240};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:472:54  */
  assign n242 = clk_gen_en[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:472:42  */
  assign n243 = {n241, n242};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:472:77  */
  assign n244 = clk_gen_en[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:472:65  */
  assign n245 = {n243, n244};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:472:100  */
  assign n246 = clk_gen_en[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:472:88  */
  assign n247 = {n245, n246};
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:482:23  */
  assign n248 = firq[15]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:483:23  */
  assign n249 = firq[7]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:484:23  */
  assign n250 = firq[14]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:485:23  */
  assign n251 = firq[13]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:486:23  */
  assign n252 = firq[12]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:487:23  */
  assign n253 = firq[11]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:488:23  */
  assign n254 = firq[10]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:489:23  */
  assign n255 = firq[8]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:490:23  */
  assign n256 = firq[5]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:491:23  */
  assign n257 = firq[6]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:492:23  */
  assign n258 = firq[2]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:493:23  */
  assign n259 = firq[9]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:494:23  */
  assign n260 = firq[4]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:495:23  */
  assign n261 = firq[3]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:496:23  */
  assign n262 = firq[1]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:497:23  */
  assign n263 = firq[0]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:505:5  */
  neorv32_cpu_0_0_4_1_40_f23860951627a2ed8cecb4a83038f47ead6bd96c core_complex_gen_n1_neorv32_cpu_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .msi_i(msw_irq),
    .mei_i(mext_irq_i),
    .mti_i(mtime_irq),
    .firq_i(cpu_firq),
    .dbi_i(dci_haltreq),
    .\icc_rx_i_icc_rx_i[rdy] (n266),
    .\icc_rx_i_icc_rx_i[ack] (n267),
    .\icc_rx_i_icc_rx_i[dat] (n268),
    .\ibus_rsp_i_ibus_rsp_i[data] (n271),
    .\ibus_rsp_i_ibus_rsp_i[ack] (n272),
    .\ibus_rsp_i_ibus_rsp_i[err] (n273),
    .\dbus_rsp_i_dbus_rsp_i[data] (n276),
    .\dbus_rsp_i_dbus_rsp_i[ack] (n277),
    .\dbus_rsp_i_dbus_rsp_i[err] (n278),
    .\icc_tx_o_icc_tx_o[rdy] (\core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[rdy] ),
    .\icc_tx_o_icc_tx_o[ack] (\core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[ack] ),
    .\icc_tx_o_icc_tx_o[dat] (\core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[dat] ),
    .\ibus_req_o_ibus_req_o[addr] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[addr] ),
    .\ibus_req_o_ibus_req_o[data] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[data] ),
    .\ibus_req_o_ibus_req_o[ben] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[ben] ),
    .\ibus_req_o_ibus_req_o[stb] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[stb] ),
    .\ibus_req_o_ibus_req_o[rw] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[rw] ),
    .\ibus_req_o_ibus_req_o[src] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[src] ),
    .\ibus_req_o_ibus_req_o[priv] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[priv] ),
    .\ibus_req_o_ibus_req_o[amo] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[amo] ),
    .\ibus_req_o_ibus_req_o[amoop] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[amoop] ),
    .\ibus_req_o_ibus_req_o[fence] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[fence] ),
    .\ibus_req_o_ibus_req_o[sleep] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[sleep] ),
    .\ibus_req_o_ibus_req_o[debug] (\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[debug] ),
    .\dbus_req_o_dbus_req_o[addr] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[addr] ),
    .\dbus_req_o_dbus_req_o[data] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[data] ),
    .\dbus_req_o_dbus_req_o[ben] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[ben] ),
    .\dbus_req_o_dbus_req_o[stb] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[stb] ),
    .\dbus_req_o_dbus_req_o[rw] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[rw] ),
    .\dbus_req_o_dbus_req_o[src] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[src] ),
    .\dbus_req_o_dbus_req_o[priv] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[priv] ),
    .\dbus_req_o_dbus_req_o[amo] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[amo] ),
    .\dbus_req_o_dbus_req_o[amoop] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[amoop] ),
    .\dbus_req_o_dbus_req_o[fence] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[fence] ),
    .\dbus_req_o_dbus_req_o[sleep] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[sleep] ),
    .\dbus_req_o_dbus_req_o[debug] (\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[debug] ));
  assign n264 = {\core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[dat] , \core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[ack] , \core_complex_gen_n1_neorv32_cpu_inst.icc_tx_o_icc_tx_o[rdy] };
  assign n266 = icc_rx[0]; // extract
  assign n267 = icc_rx[1]; // extract
  assign n268 = icc_rx[33:2]; // extract
  assign n269 = {\core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[debug] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[sleep] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[fence] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[amoop] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[amo] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[priv] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[src] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[rw] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[stb] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[ben] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[data] , \core_complex_gen_n1_neorv32_cpu_inst.ibus_req_o_ibus_req_o[addr] };
  assign n271 = cpu_i_rsp[31:0]; // extract
  assign n272 = cpu_i_rsp[32]; // extract
  assign n273 = cpu_i_rsp[33]; // extract
  assign n274 = {\core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[debug] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[sleep] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[fence] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[amoop] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[amo] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[priv] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[src] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[rw] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[stb] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[ben] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[data] , \core_complex_gen_n1_neorv32_cpu_inst.dbus_req_o_dbus_req_o[addr] };
  assign n276 = cpu_d_rsp[31:0]; // extract
  assign n277 = cpu_d_rsp[32]; // extract
  assign n278 = cpu_d_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:636:5  */
  neorv32_bus_switch_2547cc736e951fa4919853c43ae890861a3b3264 core_complex_gen_n1_neorv32_core_bus_switch_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .a_lock_i(n279),
    .\a_req_i_a_req_i[addr] (n280),
    .\a_req_i_a_req_i[data] (n281),
    .\a_req_i_a_req_i[ben] (n282),
    .\a_req_i_a_req_i[stb] (n283),
    .\a_req_i_a_req_i[rw] (n284),
    .\a_req_i_a_req_i[src] (n285),
    .\a_req_i_a_req_i[priv] (n286),
    .\a_req_i_a_req_i[amo] (n287),
    .\a_req_i_a_req_i[amoop] (n288),
    .\a_req_i_a_req_i[fence] (n289),
    .\a_req_i_a_req_i[sleep] (n290),
    .\a_req_i_a_req_i[debug] (n291),
    .\b_req_i_b_req_i[addr] (n294),
    .\b_req_i_b_req_i[data] (n295),
    .\b_req_i_b_req_i[ben] (n296),
    .\b_req_i_b_req_i[stb] (n297),
    .\b_req_i_b_req_i[rw] (n298),
    .\b_req_i_b_req_i[src] (n299),
    .\b_req_i_b_req_i[priv] (n300),
    .\b_req_i_b_req_i[amo] (n301),
    .\b_req_i_b_req_i[amoop] (n302),
    .\b_req_i_b_req_i[fence] (n303),
    .\b_req_i_b_req_i[sleep] (n304),
    .\b_req_i_b_req_i[debug] (n305),
    .\x_rsp_i_x_rsp_i[data] (n310),
    .\x_rsp_i_x_rsp_i[ack] (n311),
    .\x_rsp_i_x_rsp_i[err] (n312),
    .\a_rsp_o_a_rsp_o[data] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[data] ),
    .\a_rsp_o_a_rsp_o[ack] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[ack] ),
    .\a_rsp_o_a_rsp_o[err] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[err] ),
    .\b_rsp_o_b_rsp_o[data] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[data] ),
    .\b_rsp_o_b_rsp_o[ack] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[ack] ),
    .\b_rsp_o_b_rsp_o[err] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[err] ),
    .\x_req_o_x_req_o[addr] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[addr] ),
    .\x_req_o_x_req_o[data] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[data] ),
    .\x_req_o_x_req_o[ben] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[ben] ),
    .\x_req_o_x_req_o[stb] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[stb] ),
    .\x_req_o_x_req_o[rw] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[rw] ),
    .\x_req_o_x_req_o[src] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[src] ),
    .\x_req_o_x_req_o[priv] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[priv] ),
    .\x_req_o_x_req_o[amo] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[amo] ),
    .\x_req_o_x_req_o[amoop] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[amoop] ),
    .\x_req_o_x_req_o[fence] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[fence] ),
    .\x_req_o_x_req_o[sleep] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[sleep] ),
    .\x_req_o_x_req_o[debug] (\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[debug] ));
  assign n280 = dcache_req[31:0]; // extract
  assign n281 = dcache_req[63:32]; // extract
  assign n282 = dcache_req[67:64]; // extract
  assign n283 = dcache_req[68]; // extract
  assign n284 = dcache_req[69]; // extract
  assign n285 = dcache_req[70]; // extract
  assign n286 = dcache_req[71]; // extract
  assign n287 = dcache_req[72]; // extract
  assign n288 = dcache_req[76:73]; // extract
  assign n289 = dcache_req[77]; // extract
  assign n290 = dcache_req[78]; // extract
  assign n291 = dcache_req[79]; // extract
  assign n292 = {\core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[err] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[ack] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.a_rsp_o_a_rsp_o[data] };
  assign n294 = icache_req[31:0]; // extract
  assign n295 = icache_req[63:32]; // extract
  assign n296 = icache_req[67:64]; // extract
  assign n297 = icache_req[68]; // extract
  assign n298 = icache_req[69]; // extract
  assign n299 = icache_req[70]; // extract
  assign n300 = icache_req[71]; // extract
  assign n301 = icache_req[72]; // extract
  assign n302 = icache_req[76:73]; // extract
  assign n303 = icache_req[77]; // extract
  assign n304 = icache_req[78]; // extract
  assign n305 = icache_req[79]; // extract
  assign n306 = {\core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[err] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[ack] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.b_rsp_o_b_rsp_o[data] };
  assign n308 = {\core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[debug] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[sleep] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[fence] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[amoop] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[amo] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[priv] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[src] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[rw] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[stb] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[ben] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[data] , \core_complex_gen_n1_neorv32_core_bus_switch_inst.x_req_o_x_req_o[addr] };
  assign n310 = core_rsp[31:0]; // extract
  assign n311 = core_rsp[32]; // extract
  assign n312 = core_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:777:3  */
  neorv32_bus_gateway_15_16384_16384_268435456_2097152_d3c572afed0908e1a530126dd188e3360efa598d neorv32_bus_gateway_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\req_i_req_i[addr] (n317),
    .\req_i_req_i[data] (n318),
    .\req_i_req_i[ben] (n319),
    .\req_i_req_i[stb] (n320),
    .\req_i_req_i[rw] (n321),
    .\req_i_req_i[src] (n322),
    .\req_i_req_i[priv] (n323),
    .\req_i_req_i[amo] (n324),
    .\req_i_req_i[amoop] (n325),
    .\req_i_req_i[fence] (n326),
    .\req_i_req_i[sleep] (n327),
    .\req_i_req_i[debug] (n328),
    .\a_rsp_i_a_rsp_i[data] (n333),
    .\a_rsp_i_a_rsp_i[ack] (n334),
    .\a_rsp_i_a_rsp_i[err] (n335),
    .\b_rsp_i_b_rsp_i[data] (n338),
    .\b_rsp_i_b_rsp_i[ack] (n339),
    .\b_rsp_i_b_rsp_i[err] (n340),
    .\c_rsp_i_c_rsp_i[data] (n343),
    .\c_rsp_i_c_rsp_i[ack] (n344),
    .\c_rsp_i_c_rsp_i[err] (n345),
    .\d_rsp_i_d_rsp_i[data] (n348),
    .\d_rsp_i_d_rsp_i[ack] (n349),
    .\d_rsp_i_d_rsp_i[err] (n350),
    .\x_rsp_i_x_rsp_i[data] (n353),
    .\x_rsp_i_x_rsp_i[ack] (n354),
    .\x_rsp_i_x_rsp_i[err] (n355),
    .\rsp_o_rsp_o[data] (\neorv32_bus_gateway_inst.rsp_o_rsp_o[data] ),
    .\rsp_o_rsp_o[ack] (\neorv32_bus_gateway_inst.rsp_o_rsp_o[ack] ),
    .\rsp_o_rsp_o[err] (\neorv32_bus_gateway_inst.rsp_o_rsp_o[err] ),
    .\a_req_o_a_req_o[addr] (),
    .\a_req_o_a_req_o[data] (),
    .\a_req_o_a_req_o[ben] (),
    .\a_req_o_a_req_o[stb] (),
    .\a_req_o_a_req_o[rw] (),
    .\a_req_o_a_req_o[src] (),
    .\a_req_o_a_req_o[priv] (),
    .\a_req_o_a_req_o[amo] (),
    .\a_req_o_a_req_o[amoop] (),
    .\a_req_o_a_req_o[fence] (),
    .\a_req_o_a_req_o[sleep] (),
    .\a_req_o_a_req_o[debug] (),
    .\b_req_o_b_req_o[addr] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[addr] ),
    .\b_req_o_b_req_o[data] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[data] ),
    .\b_req_o_b_req_o[ben] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[ben] ),
    .\b_req_o_b_req_o[stb] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[stb] ),
    .\b_req_o_b_req_o[rw] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[rw] ),
    .\b_req_o_b_req_o[src] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[src] ),
    .\b_req_o_b_req_o[priv] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[priv] ),
    .\b_req_o_b_req_o[amo] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[amo] ),
    .\b_req_o_b_req_o[amoop] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[amoop] ),
    .\b_req_o_b_req_o[fence] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[fence] ),
    .\b_req_o_b_req_o[sleep] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[sleep] ),
    .\b_req_o_b_req_o[debug] (\neorv32_bus_gateway_inst.b_req_o_b_req_o[debug] ),
    .\c_req_o_c_req_o[addr] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[addr] ),
    .\c_req_o_c_req_o[data] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[data] ),
    .\c_req_o_c_req_o[ben] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[ben] ),
    .\c_req_o_c_req_o[stb] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[stb] ),
    .\c_req_o_c_req_o[rw] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[rw] ),
    .\c_req_o_c_req_o[src] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[src] ),
    .\c_req_o_c_req_o[priv] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[priv] ),
    .\c_req_o_c_req_o[amo] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[amo] ),
    .\c_req_o_c_req_o[amoop] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[amoop] ),
    .\c_req_o_c_req_o[fence] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[fence] ),
    .\c_req_o_c_req_o[sleep] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[sleep] ),
    .\c_req_o_c_req_o[debug] (\neorv32_bus_gateway_inst.c_req_o_c_req_o[debug] ),
    .\d_req_o_d_req_o[addr] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[addr] ),
    .\d_req_o_d_req_o[data] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[data] ),
    .\d_req_o_d_req_o[ben] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[ben] ),
    .\d_req_o_d_req_o[stb] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[stb] ),
    .\d_req_o_d_req_o[rw] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[rw] ),
    .\d_req_o_d_req_o[src] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[src] ),
    .\d_req_o_d_req_o[priv] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[priv] ),
    .\d_req_o_d_req_o[amo] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[amo] ),
    .\d_req_o_d_req_o[amoop] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[amoop] ),
    .\d_req_o_d_req_o[fence] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[fence] ),
    .\d_req_o_d_req_o[sleep] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[sleep] ),
    .\d_req_o_d_req_o[debug] (\neorv32_bus_gateway_inst.d_req_o_d_req_o[debug] ),
    .\x_req_o_x_req_o[addr] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[addr] ),
    .\x_req_o_x_req_o[data] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[data] ),
    .\x_req_o_x_req_o[ben] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[ben] ),
    .\x_req_o_x_req_o[stb] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[stb] ),
    .\x_req_o_x_req_o[rw] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[rw] ),
    .\x_req_o_x_req_o[src] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[src] ),
    .\x_req_o_x_req_o[priv] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[priv] ),
    .\x_req_o_x_req_o[amo] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[amo] ),
    .\x_req_o_x_req_o[amoop] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[amoop] ),
    .\x_req_o_x_req_o[fence] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[fence] ),
    .\x_req_o_x_req_o[sleep] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[sleep] ),
    .\x_req_o_x_req_o[debug] (\neorv32_bus_gateway_inst.x_req_o_x_req_o[debug] ));
  assign n317 = sys3_req[31:0]; // extract
  assign n318 = sys3_req[63:32]; // extract
  assign n319 = sys3_req[67:64]; // extract
  assign n320 = sys3_req[68]; // extract
  assign n321 = sys3_req[69]; // extract
  assign n322 = sys3_req[70]; // extract
  assign n323 = sys3_req[71]; // extract
  assign n324 = sys3_req[72]; // extract
  assign n325 = sys3_req[76:73]; // extract
  assign n326 = sys3_req[77]; // extract
  assign n327 = sys3_req[78]; // extract
  assign n328 = sys3_req[79]; // extract
  assign n329 = {\neorv32_bus_gateway_inst.rsp_o_rsp_o[err] , \neorv32_bus_gateway_inst.rsp_o_rsp_o[ack] , \neorv32_bus_gateway_inst.rsp_o_rsp_o[data] };
  assign n333 = imem_rsp[31:0]; // extract
  assign n334 = imem_rsp[32]; // extract
  assign n335 = imem_rsp[33]; // extract
  assign n336 = {\neorv32_bus_gateway_inst.b_req_o_b_req_o[debug] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[sleep] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[fence] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[amoop] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[amo] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[priv] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[src] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[rw] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[stb] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[ben] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[data] , \neorv32_bus_gateway_inst.b_req_o_b_req_o[addr] };
  assign n338 = dmem_rsp[31:0]; // extract
  assign n339 = dmem_rsp[32]; // extract
  assign n340 = dmem_rsp[33]; // extract
  assign n341 = {\neorv32_bus_gateway_inst.c_req_o_c_req_o[debug] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[sleep] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[fence] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[amoop] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[amo] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[priv] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[src] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[rw] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[stb] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[ben] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[data] , \neorv32_bus_gateway_inst.c_req_o_c_req_o[addr] };
  assign n343 = xip_rsp[31:0]; // extract
  assign n344 = xip_rsp[32]; // extract
  assign n345 = xip_rsp[33]; // extract
  assign n346 = {\neorv32_bus_gateway_inst.d_req_o_d_req_o[debug] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[sleep] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[fence] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[amoop] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[amo] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[priv] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[src] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[rw] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[stb] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[ben] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[data] , \neorv32_bus_gateway_inst.d_req_o_d_req_o[addr] };
  assign n348 = io_rsp[31:0]; // extract
  assign n349 = io_rsp[32]; // extract
  assign n350 = io_rsp[33]; // extract
  assign n351 = {\neorv32_bus_gateway_inst.x_req_o_x_req_o[debug] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[sleep] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[fence] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[amoop] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[amo] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[priv] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[src] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[rw] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[stb] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[ben] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[data] , \neorv32_bus_gateway_inst.x_req_o_x_req_o[addr] };
  assign n353 = xbus_rsp[31:0]; // extract
  assign n354 = xbus_rsp[32]; // extract
  assign n355 = xbus_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:859:7  */
  neorv32_dmem_16384 memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n357),
    .\bus_req_i_bus_req_i[data] (n358),
    .\bus_req_i_bus_req_i[ben] (n359),
    .\bus_req_i_bus_req_i[stb] (n360),
    .\bus_req_i_bus_req_i[rw] (n361),
    .\bus_req_i_bus_req_i[src] (n362),
    .\bus_req_i_bus_req_i[priv] (n363),
    .\bus_req_i_bus_req_i[amo] (n364),
    .\bus_req_i_bus_req_i[amoop] (n365),
    .\bus_req_i_bus_req_i[fence] (n366),
    .\bus_req_i_bus_req_i[sleep] (n367),
    .\bus_req_i_bus_req_i[debug] (n368),
    .\bus_rsp_o_bus_rsp_o[data] (\memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[err] ));
  assign n357 = dmem_req[31:0]; // extract
  assign n358 = dmem_req[63:32]; // extract
  assign n359 = dmem_req[67:64]; // extract
  assign n360 = dmem_req[68]; // extract
  assign n361 = dmem_req[69]; // extract
  assign n362 = dmem_req[70]; // extract
  assign n363 = dmem_req[71]; // extract
  assign n364 = dmem_req[72]; // extract
  assign n365 = dmem_req[76:73]; // extract
  assign n366 = dmem_req[77]; // extract
  assign n367 = dmem_req[78]; // extract
  assign n368 = dmem_req[79]; // extract
  assign n369 = {\memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[err] , \memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[ack] , \memory_system_neorv32_int_dmem_enabled_neorv32_int_dmem_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:883:7  */
  neorv32_xip_bf8b4530d8d246dd74ac53a13471bba17941dff7 memory_system_neorv32_xip_enabled_neorv32_xip_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n372),
    .\bus_req_i_bus_req_i[data] (n373),
    .\bus_req_i_bus_req_i[ben] (n374),
    .\bus_req_i_bus_req_i[stb] (n375),
    .\bus_req_i_bus_req_i[rw] (n376),
    .\bus_req_i_bus_req_i[src] (n377),
    .\bus_req_i_bus_req_i[priv] (n378),
    .\bus_req_i_bus_req_i[amo] (n379),
    .\bus_req_i_bus_req_i[amoop] (n380),
    .\bus_req_i_bus_req_i[fence] (n381),
    .\bus_req_i_bus_req_i[sleep] (n382),
    .\bus_req_i_bus_req_i[debug] (n383),
    .\xip_req_i_xip_req_i[addr] (n386),
    .\xip_req_i_xip_req_i[data] (n387),
    .\xip_req_i_xip_req_i[ben] (n388),
    .\xip_req_i_xip_req_i[stb] (n389),
    .\xip_req_i_xip_req_i[rw] (n390),
    .\xip_req_i_xip_req_i[src] (n391),
    .\xip_req_i_xip_req_i[priv] (n392),
    .\xip_req_i_xip_req_i[amo] (n393),
    .\xip_req_i_xip_req_i[amoop] (n394),
    .\xip_req_i_xip_req_i[fence] (n395),
    .\xip_req_i_xip_req_i[sleep] (n396),
    .\xip_req_i_xip_req_i[debug] (n397),
    .clkgen_i(clk_gen),
    .spi_dat_i(xip_dat_i),
    .\bus_rsp_o_bus_rsp_o[data] (\memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[err] ),
    .\xip_rsp_o_xip_rsp_o[data] (\memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[data] ),
    .\xip_rsp_o_xip_rsp_o[ack] (\memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[ack] ),
    .\xip_rsp_o_xip_rsp_o[err] (\memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[err] ),
    .clkgen_en_o(\memory_system_neorv32_xip_enabled_neorv32_xip_inst.clkgen_en_o ),
    .spi_csn_o(\memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_csn_o ),
    .spi_clk_o(\memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_clk_o ),
    .spi_dat_o(\memory_system_neorv32_xip_enabled_neorv32_xip_inst.spi_dat_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:890:33  */
  assign n371 = iodev_req[479:400]; // extract
  assign n372 = n371[31:0]; // extract
  assign n373 = n371[63:32]; // extract
  assign n374 = n371[67:64]; // extract
  assign n375 = n371[68]; // extract
  assign n376 = n371[69]; // extract
  assign n377 = n371[70]; // extract
  assign n378 = n371[71]; // extract
  assign n379 = n371[72]; // extract
  assign n380 = n371[76:73]; // extract
  assign n381 = n371[77]; // extract
  assign n382 = n371[78]; // extract
  assign n383 = n371[79]; // extract
  assign n384 = {\memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[err] , \memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[ack] , \memory_system_neorv32_xip_enabled_neorv32_xip_inst.bus_rsp_o_bus_rsp_o[data] };
  assign n386 = xipcache_req[31:0]; // extract
  assign n387 = xipcache_req[63:32]; // extract
  assign n388 = xipcache_req[67:64]; // extract
  assign n389 = xipcache_req[68]; // extract
  assign n390 = xipcache_req[69]; // extract
  assign n391 = xipcache_req[70]; // extract
  assign n392 = xipcache_req[71]; // extract
  assign n393 = xipcache_req[72]; // extract
  assign n394 = xipcache_req[76:73]; // extract
  assign n395 = xipcache_req[77]; // extract
  assign n396 = xipcache_req[78]; // extract
  assign n397 = xipcache_req[79]; // extract
  assign n398 = {\memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[err] , \memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[ack] , \memory_system_neorv32_xip_enabled_neorv32_xip_inst.xip_rsp_o_xip_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:905:9  */
  neorv32_cache_16_64_69f24bf1e9d58f38577f662be0ab41a8f51212bb memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\host_req_i_host_req_i[addr] (n404),
    .\host_req_i_host_req_i[data] (n405),
    .\host_req_i_host_req_i[ben] (n406),
    .\host_req_i_host_req_i[stb] (n407),
    .\host_req_i_host_req_i[rw] (n408),
    .\host_req_i_host_req_i[src] (n409),
    .\host_req_i_host_req_i[priv] (n410),
    .\host_req_i_host_req_i[amo] (n411),
    .\host_req_i_host_req_i[amoop] (n412),
    .\host_req_i_host_req_i[fence] (n413),
    .\host_req_i_host_req_i[sleep] (n414),
    .\host_req_i_host_req_i[debug] (n415),
    .\bus_rsp_i_bus_rsp_i[data] (n420),
    .\bus_rsp_i_bus_rsp_i[ack] (n421),
    .\bus_rsp_i_bus_rsp_i[err] (n422),
    .\host_rsp_o_host_rsp_o[data] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[data] ),
    .\host_rsp_o_host_rsp_o[ack] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[ack] ),
    .\host_rsp_o_host_rsp_o[err] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[err] ),
    .\bus_req_o_bus_req_o[addr] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[addr] ),
    .\bus_req_o_bus_req_o[data] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[data] ),
    .\bus_req_o_bus_req_o[ben] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[ben] ),
    .\bus_req_o_bus_req_o[stb] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[stb] ),
    .\bus_req_o_bus_req_o[rw] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[rw] ),
    .\bus_req_o_bus_req_o[src] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[src] ),
    .\bus_req_o_bus_req_o[priv] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[priv] ),
    .\bus_req_o_bus_req_o[amo] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[amo] ),
    .\bus_req_o_bus_req_o[amoop] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[amoop] ),
    .\bus_req_o_bus_req_o[fence] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[fence] ),
    .\bus_req_o_bus_req_o[sleep] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[sleep] ),
    .\bus_req_o_bus_req_o[debug] (\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[debug] ));
  assign n404 = xip_req[31:0]; // extract
  assign n405 = xip_req[63:32]; // extract
  assign n406 = xip_req[67:64]; // extract
  assign n407 = xip_req[68]; // extract
  assign n408 = xip_req[69]; // extract
  assign n409 = xip_req[70]; // extract
  assign n410 = xip_req[71]; // extract
  assign n411 = xip_req[72]; // extract
  assign n412 = xip_req[76:73]; // extract
  assign n413 = xip_req[77]; // extract
  assign n414 = xip_req[78]; // extract
  assign n415 = xip_req[79]; // extract
  assign n416 = {\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[err] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[ack] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.host_rsp_o_host_rsp_o[data] };
  assign n418 = {\memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[debug] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[sleep] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[fence] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[amoop] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[amo] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[priv] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[src] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[rw] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[stb] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[ben] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[data] , \memory_system_neorv32_xip_enabled_neorv32_xipcache_enabled_neorv32_xcache_inst.bus_req_o_bus_req_o[addr] };
  assign n420 = xipcache_rsp[31:0]; // extract
  assign n421 = xipcache_rsp[32]; // extract
  assign n422 = xipcache_rsp[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:948:7  */
  neorv32_xbus_255_5ba93c9db0cff93f52b521d7420e43f6eda2784f memory_system_neorv32_xbus_enabled_neorv32_xbus_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n423),
    .\bus_req_i_bus_req_i[data] (n424),
    .\bus_req_i_bus_req_i[ben] (n425),
    .\bus_req_i_bus_req_i[stb] (n426),
    .\bus_req_i_bus_req_i[rw] (n427),
    .\bus_req_i_bus_req_i[src] (n428),
    .\bus_req_i_bus_req_i[priv] (n429),
    .\bus_req_i_bus_req_i[amo] (n430),
    .\bus_req_i_bus_req_i[amoop] (n431),
    .\bus_req_i_bus_req_i[fence] (n432),
    .\bus_req_i_bus_req_i[sleep] (n433),
    .\bus_req_i_bus_req_i[debug] (n434),
    .xbus_dat_i(xbus_dat_i),
    .xbus_ack_i(xbus_ack_i),
    .xbus_err_i(xbus_err_i),
    .\bus_rsp_o_bus_rsp_o[data] (\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[err] ),
    .xbus_adr_o(\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_adr_o ),
    .xbus_dat_o(\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_dat_o ),
    .xbus_tag_o(\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_tag_o ),
    .xbus_we_o(\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_we_o ),
    .xbus_sel_o(\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_sel_o ),
    .xbus_stb_o(\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_stb_o ),
    .xbus_cyc_o(\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.xbus_cyc_o ));
  assign n423 = xcache_req[31:0]; // extract
  assign n424 = xcache_req[63:32]; // extract
  assign n425 = xcache_req[67:64]; // extract
  assign n426 = xcache_req[68]; // extract
  assign n427 = xcache_req[69]; // extract
  assign n428 = xcache_req[70]; // extract
  assign n429 = xcache_req[71]; // extract
  assign n430 = xcache_req[72]; // extract
  assign n431 = xcache_req[76:73]; // extract
  assign n432 = xcache_req[77]; // extract
  assign n433 = xcache_req[78]; // extract
  assign n434 = xcache_req[79]; // extract
  assign n435 = {\memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[err] , \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[ack] , \memory_system_neorv32_xbus_enabled_neorv32_xbus_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1024:5  */
  neorv32_bus_io_switch_65536_19a0518872770ca4a65ad41d181dd3070f957778 io_system_neorv32_bus_io_switch_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\main_req_i_main_req_i[addr] (n444),
    .\main_req_i_main_req_i[data] (n445),
    .\main_req_i_main_req_i[ben] (n446),
    .\main_req_i_main_req_i[stb] (n447),
    .\main_req_i_main_req_i[rw] (n448),
    .\main_req_i_main_req_i[src] (n449),
    .\main_req_i_main_req_i[priv] (n450),
    .\main_req_i_main_req_i[amo] (n451),
    .\main_req_i_main_req_i[amoop] (n452),
    .\main_req_i_main_req_i[fence] (n453),
    .\main_req_i_main_req_i[sleep] (n454),
    .\main_req_i_main_req_i[debug] (n455),
    .\dev_00_rsp_i_dev_00_rsp_i[data] (n461),
    .\dev_00_rsp_i_dev_00_rsp_i[ack] (n462),
    .\dev_00_rsp_i_dev_00_rsp_i[err] (n463),
    .\dev_01_rsp_i_dev_01_rsp_i[data] (n465),
    .\dev_01_rsp_i_dev_01_rsp_i[ack] (n466),
    .\dev_01_rsp_i_dev_01_rsp_i[err] (n467),
    .\dev_02_rsp_i_dev_02_rsp_i[data] (n469),
    .\dev_02_rsp_i_dev_02_rsp_i[ack] (n470),
    .\dev_02_rsp_i_dev_02_rsp_i[err] (n471),
    .\dev_03_rsp_i_dev_03_rsp_i[data] (n473),
    .\dev_03_rsp_i_dev_03_rsp_i[ack] (n474),
    .\dev_03_rsp_i_dev_03_rsp_i[err] (n475),
    .\dev_04_rsp_i_dev_04_rsp_i[data] (n477),
    .\dev_04_rsp_i_dev_04_rsp_i[ack] (n478),
    .\dev_04_rsp_i_dev_04_rsp_i[err] (n479),
    .\dev_05_rsp_i_dev_05_rsp_i[data] (n481),
    .\dev_05_rsp_i_dev_05_rsp_i[ack] (n482),
    .\dev_05_rsp_i_dev_05_rsp_i[err] (n483),
    .\dev_06_rsp_i_dev_06_rsp_i[data] (n485),
    .\dev_06_rsp_i_dev_06_rsp_i[ack] (n486),
    .\dev_06_rsp_i_dev_06_rsp_i[err] (n487),
    .\dev_07_rsp_i_dev_07_rsp_i[data] (n489),
    .\dev_07_rsp_i_dev_07_rsp_i[ack] (n490),
    .\dev_07_rsp_i_dev_07_rsp_i[err] (n491),
    .\dev_08_rsp_i_dev_08_rsp_i[data] (n493),
    .\dev_08_rsp_i_dev_08_rsp_i[ack] (n494),
    .\dev_08_rsp_i_dev_08_rsp_i[err] (n495),
    .\dev_09_rsp_i_dev_09_rsp_i[data] (n497),
    .\dev_09_rsp_i_dev_09_rsp_i[ack] (n498),
    .\dev_09_rsp_i_dev_09_rsp_i[err] (n499),
    .\dev_10_rsp_i_dev_10_rsp_i[data] (n503),
    .\dev_10_rsp_i_dev_10_rsp_i[ack] (n504),
    .\dev_10_rsp_i_dev_10_rsp_i[err] (n505),
    .\dev_11_rsp_i_dev_11_rsp_i[data] (n509),
    .\dev_11_rsp_i_dev_11_rsp_i[ack] (n510),
    .\dev_11_rsp_i_dev_11_rsp_i[err] (n511),
    .\dev_12_rsp_i_dev_12_rsp_i[data] (n515),
    .\dev_12_rsp_i_dev_12_rsp_i[ack] (n516),
    .\dev_12_rsp_i_dev_12_rsp_i[err] (n517),
    .\dev_13_rsp_i_dev_13_rsp_i[data] (n521),
    .\dev_13_rsp_i_dev_13_rsp_i[ack] (n522),
    .\dev_13_rsp_i_dev_13_rsp_i[err] (n523),
    .\dev_14_rsp_i_dev_14_rsp_i[data] (n527),
    .\dev_14_rsp_i_dev_14_rsp_i[ack] (n528),
    .\dev_14_rsp_i_dev_14_rsp_i[err] (n529),
    .\dev_15_rsp_i_dev_15_rsp_i[data] (n533),
    .\dev_15_rsp_i_dev_15_rsp_i[ack] (n534),
    .\dev_15_rsp_i_dev_15_rsp_i[err] (n535),
    .\dev_16_rsp_i_dev_16_rsp_i[data] (n539),
    .\dev_16_rsp_i_dev_16_rsp_i[ack] (n540),
    .\dev_16_rsp_i_dev_16_rsp_i[err] (n541),
    .\dev_17_rsp_i_dev_17_rsp_i[data] (n545),
    .\dev_17_rsp_i_dev_17_rsp_i[ack] (n546),
    .\dev_17_rsp_i_dev_17_rsp_i[err] (n547),
    .\dev_18_rsp_i_dev_18_rsp_i[data] (n551),
    .\dev_18_rsp_i_dev_18_rsp_i[ack] (n552),
    .\dev_18_rsp_i_dev_18_rsp_i[err] (n553),
    .\dev_19_rsp_i_dev_19_rsp_i[data] (n555),
    .\dev_19_rsp_i_dev_19_rsp_i[ack] (n556),
    .\dev_19_rsp_i_dev_19_rsp_i[err] (n557),
    .\dev_20_rsp_i_dev_20_rsp_i[data] (n561),
    .\dev_20_rsp_i_dev_20_rsp_i[ack] (n562),
    .\dev_20_rsp_i_dev_20_rsp_i[err] (n563),
    .\dev_21_rsp_i_dev_21_rsp_i[data] (n567),
    .\dev_21_rsp_i_dev_21_rsp_i[ack] (n568),
    .\dev_21_rsp_i_dev_21_rsp_i[err] (n569),
    .\dev_22_rsp_i_dev_22_rsp_i[data] (n573),
    .\dev_22_rsp_i_dev_22_rsp_i[ack] (n574),
    .\dev_22_rsp_i_dev_22_rsp_i[err] (n575),
    .\dev_23_rsp_i_dev_23_rsp_i[data] (n579),
    .\dev_23_rsp_i_dev_23_rsp_i[ack] (n580),
    .\dev_23_rsp_i_dev_23_rsp_i[err] (n581),
    .\dev_24_rsp_i_dev_24_rsp_i[data] (n585),
    .\dev_24_rsp_i_dev_24_rsp_i[ack] (n586),
    .\dev_24_rsp_i_dev_24_rsp_i[err] (n587),
    .\dev_25_rsp_i_dev_25_rsp_i[data] (n591),
    .\dev_25_rsp_i_dev_25_rsp_i[ack] (n592),
    .\dev_25_rsp_i_dev_25_rsp_i[err] (n593),
    .\dev_26_rsp_i_dev_26_rsp_i[data] (n597),
    .\dev_26_rsp_i_dev_26_rsp_i[ack] (n598),
    .\dev_26_rsp_i_dev_26_rsp_i[err] (n599),
    .\dev_27_rsp_i_dev_27_rsp_i[data] (n603),
    .\dev_27_rsp_i_dev_27_rsp_i[ack] (n604),
    .\dev_27_rsp_i_dev_27_rsp_i[err] (n605),
    .\dev_28_rsp_i_dev_28_rsp_i[data] (n609),
    .\dev_28_rsp_i_dev_28_rsp_i[ack] (n610),
    .\dev_28_rsp_i_dev_28_rsp_i[err] (n611),
    .\dev_29_rsp_i_dev_29_rsp_i[data] (n615),
    .\dev_29_rsp_i_dev_29_rsp_i[ack] (n616),
    .\dev_29_rsp_i_dev_29_rsp_i[err] (n617),
    .\dev_30_rsp_i_dev_30_rsp_i[data] (n621),
    .\dev_30_rsp_i_dev_30_rsp_i[ack] (n622),
    .\dev_30_rsp_i_dev_30_rsp_i[err] (n623),
    .\dev_31_rsp_i_dev_31_rsp_i[data] (n627),
    .\dev_31_rsp_i_dev_31_rsp_i[ack] (n628),
    .\dev_31_rsp_i_dev_31_rsp_i[err] (n629),
    .\main_rsp_o_main_rsp_o[data] (\io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[data] ),
    .\main_rsp_o_main_rsp_o[ack] (\io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[ack] ),
    .\main_rsp_o_main_rsp_o[err] (\io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[err] ),
    .\dev_00_req_o_dev_00_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[addr] ),
    .\dev_00_req_o_dev_00_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[data] ),
    .\dev_00_req_o_dev_00_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[ben] ),
    .\dev_00_req_o_dev_00_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[stb] ),
    .\dev_00_req_o_dev_00_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[rw] ),
    .\dev_00_req_o_dev_00_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[src] ),
    .\dev_00_req_o_dev_00_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[priv] ),
    .\dev_00_req_o_dev_00_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[amo] ),
    .\dev_00_req_o_dev_00_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[amoop] ),
    .\dev_00_req_o_dev_00_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[fence] ),
    .\dev_00_req_o_dev_00_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[sleep] ),
    .\dev_00_req_o_dev_00_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[debug] ),
    .\dev_01_req_o_dev_01_req_o[addr] (),
    .\dev_01_req_o_dev_01_req_o[data] (),
    .\dev_01_req_o_dev_01_req_o[ben] (),
    .\dev_01_req_o_dev_01_req_o[stb] (),
    .\dev_01_req_o_dev_01_req_o[rw] (),
    .\dev_01_req_o_dev_01_req_o[src] (),
    .\dev_01_req_o_dev_01_req_o[priv] (),
    .\dev_01_req_o_dev_01_req_o[amo] (),
    .\dev_01_req_o_dev_01_req_o[amoop] (),
    .\dev_01_req_o_dev_01_req_o[fence] (),
    .\dev_01_req_o_dev_01_req_o[sleep] (),
    .\dev_01_req_o_dev_01_req_o[debug] (),
    .\dev_02_req_o_dev_02_req_o[addr] (),
    .\dev_02_req_o_dev_02_req_o[data] (),
    .\dev_02_req_o_dev_02_req_o[ben] (),
    .\dev_02_req_o_dev_02_req_o[stb] (),
    .\dev_02_req_o_dev_02_req_o[rw] (),
    .\dev_02_req_o_dev_02_req_o[src] (),
    .\dev_02_req_o_dev_02_req_o[priv] (),
    .\dev_02_req_o_dev_02_req_o[amo] (),
    .\dev_02_req_o_dev_02_req_o[amoop] (),
    .\dev_02_req_o_dev_02_req_o[fence] (),
    .\dev_02_req_o_dev_02_req_o[sleep] (),
    .\dev_02_req_o_dev_02_req_o[debug] (),
    .\dev_03_req_o_dev_03_req_o[addr] (),
    .\dev_03_req_o_dev_03_req_o[data] (),
    .\dev_03_req_o_dev_03_req_o[ben] (),
    .\dev_03_req_o_dev_03_req_o[stb] (),
    .\dev_03_req_o_dev_03_req_o[rw] (),
    .\dev_03_req_o_dev_03_req_o[src] (),
    .\dev_03_req_o_dev_03_req_o[priv] (),
    .\dev_03_req_o_dev_03_req_o[amo] (),
    .\dev_03_req_o_dev_03_req_o[amoop] (),
    .\dev_03_req_o_dev_03_req_o[fence] (),
    .\dev_03_req_o_dev_03_req_o[sleep] (),
    .\dev_03_req_o_dev_03_req_o[debug] (),
    .\dev_04_req_o_dev_04_req_o[addr] (),
    .\dev_04_req_o_dev_04_req_o[data] (),
    .\dev_04_req_o_dev_04_req_o[ben] (),
    .\dev_04_req_o_dev_04_req_o[stb] (),
    .\dev_04_req_o_dev_04_req_o[rw] (),
    .\dev_04_req_o_dev_04_req_o[src] (),
    .\dev_04_req_o_dev_04_req_o[priv] (),
    .\dev_04_req_o_dev_04_req_o[amo] (),
    .\dev_04_req_o_dev_04_req_o[amoop] (),
    .\dev_04_req_o_dev_04_req_o[fence] (),
    .\dev_04_req_o_dev_04_req_o[sleep] (),
    .\dev_04_req_o_dev_04_req_o[debug] (),
    .\dev_05_req_o_dev_05_req_o[addr] (),
    .\dev_05_req_o_dev_05_req_o[data] (),
    .\dev_05_req_o_dev_05_req_o[ben] (),
    .\dev_05_req_o_dev_05_req_o[stb] (),
    .\dev_05_req_o_dev_05_req_o[rw] (),
    .\dev_05_req_o_dev_05_req_o[src] (),
    .\dev_05_req_o_dev_05_req_o[priv] (),
    .\dev_05_req_o_dev_05_req_o[amo] (),
    .\dev_05_req_o_dev_05_req_o[amoop] (),
    .\dev_05_req_o_dev_05_req_o[fence] (),
    .\dev_05_req_o_dev_05_req_o[sleep] (),
    .\dev_05_req_o_dev_05_req_o[debug] (),
    .\dev_06_req_o_dev_06_req_o[addr] (),
    .\dev_06_req_o_dev_06_req_o[data] (),
    .\dev_06_req_o_dev_06_req_o[ben] (),
    .\dev_06_req_o_dev_06_req_o[stb] (),
    .\dev_06_req_o_dev_06_req_o[rw] (),
    .\dev_06_req_o_dev_06_req_o[src] (),
    .\dev_06_req_o_dev_06_req_o[priv] (),
    .\dev_06_req_o_dev_06_req_o[amo] (),
    .\dev_06_req_o_dev_06_req_o[amoop] (),
    .\dev_06_req_o_dev_06_req_o[fence] (),
    .\dev_06_req_o_dev_06_req_o[sleep] (),
    .\dev_06_req_o_dev_06_req_o[debug] (),
    .\dev_07_req_o_dev_07_req_o[addr] (),
    .\dev_07_req_o_dev_07_req_o[data] (),
    .\dev_07_req_o_dev_07_req_o[ben] (),
    .\dev_07_req_o_dev_07_req_o[stb] (),
    .\dev_07_req_o_dev_07_req_o[rw] (),
    .\dev_07_req_o_dev_07_req_o[src] (),
    .\dev_07_req_o_dev_07_req_o[priv] (),
    .\dev_07_req_o_dev_07_req_o[amo] (),
    .\dev_07_req_o_dev_07_req_o[amoop] (),
    .\dev_07_req_o_dev_07_req_o[fence] (),
    .\dev_07_req_o_dev_07_req_o[sleep] (),
    .\dev_07_req_o_dev_07_req_o[debug] (),
    .\dev_08_req_o_dev_08_req_o[addr] (),
    .\dev_08_req_o_dev_08_req_o[data] (),
    .\dev_08_req_o_dev_08_req_o[ben] (),
    .\dev_08_req_o_dev_08_req_o[stb] (),
    .\dev_08_req_o_dev_08_req_o[rw] (),
    .\dev_08_req_o_dev_08_req_o[src] (),
    .\dev_08_req_o_dev_08_req_o[priv] (),
    .\dev_08_req_o_dev_08_req_o[amo] (),
    .\dev_08_req_o_dev_08_req_o[amoop] (),
    .\dev_08_req_o_dev_08_req_o[fence] (),
    .\dev_08_req_o_dev_08_req_o[sleep] (),
    .\dev_08_req_o_dev_08_req_o[debug] (),
    .\dev_09_req_o_dev_09_req_o[addr] (),
    .\dev_09_req_o_dev_09_req_o[data] (),
    .\dev_09_req_o_dev_09_req_o[ben] (),
    .\dev_09_req_o_dev_09_req_o[stb] (),
    .\dev_09_req_o_dev_09_req_o[rw] (),
    .\dev_09_req_o_dev_09_req_o[src] (),
    .\dev_09_req_o_dev_09_req_o[priv] (),
    .\dev_09_req_o_dev_09_req_o[amo] (),
    .\dev_09_req_o_dev_09_req_o[amoop] (),
    .\dev_09_req_o_dev_09_req_o[fence] (),
    .\dev_09_req_o_dev_09_req_o[sleep] (),
    .\dev_09_req_o_dev_09_req_o[debug] (),
    .\dev_10_req_o_dev_10_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[addr] ),
    .\dev_10_req_o_dev_10_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[data] ),
    .\dev_10_req_o_dev_10_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[ben] ),
    .\dev_10_req_o_dev_10_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[stb] ),
    .\dev_10_req_o_dev_10_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[rw] ),
    .\dev_10_req_o_dev_10_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[src] ),
    .\dev_10_req_o_dev_10_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[priv] ),
    .\dev_10_req_o_dev_10_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[amo] ),
    .\dev_10_req_o_dev_10_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[amoop] ),
    .\dev_10_req_o_dev_10_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[fence] ),
    .\dev_10_req_o_dev_10_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[sleep] ),
    .\dev_10_req_o_dev_10_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[debug] ),
    .\dev_11_req_o_dev_11_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[addr] ),
    .\dev_11_req_o_dev_11_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[data] ),
    .\dev_11_req_o_dev_11_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[ben] ),
    .\dev_11_req_o_dev_11_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[stb] ),
    .\dev_11_req_o_dev_11_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[rw] ),
    .\dev_11_req_o_dev_11_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[src] ),
    .\dev_11_req_o_dev_11_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[priv] ),
    .\dev_11_req_o_dev_11_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[amo] ),
    .\dev_11_req_o_dev_11_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[amoop] ),
    .\dev_11_req_o_dev_11_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[fence] ),
    .\dev_11_req_o_dev_11_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[sleep] ),
    .\dev_11_req_o_dev_11_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[debug] ),
    .\dev_12_req_o_dev_12_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[addr] ),
    .\dev_12_req_o_dev_12_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[data] ),
    .\dev_12_req_o_dev_12_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[ben] ),
    .\dev_12_req_o_dev_12_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[stb] ),
    .\dev_12_req_o_dev_12_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[rw] ),
    .\dev_12_req_o_dev_12_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[src] ),
    .\dev_12_req_o_dev_12_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[priv] ),
    .\dev_12_req_o_dev_12_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[amo] ),
    .\dev_12_req_o_dev_12_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[amoop] ),
    .\dev_12_req_o_dev_12_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[fence] ),
    .\dev_12_req_o_dev_12_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[sleep] ),
    .\dev_12_req_o_dev_12_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[debug] ),
    .\dev_13_req_o_dev_13_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[addr] ),
    .\dev_13_req_o_dev_13_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[data] ),
    .\dev_13_req_o_dev_13_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[ben] ),
    .\dev_13_req_o_dev_13_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[stb] ),
    .\dev_13_req_o_dev_13_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[rw] ),
    .\dev_13_req_o_dev_13_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[src] ),
    .\dev_13_req_o_dev_13_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[priv] ),
    .\dev_13_req_o_dev_13_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[amo] ),
    .\dev_13_req_o_dev_13_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[amoop] ),
    .\dev_13_req_o_dev_13_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[fence] ),
    .\dev_13_req_o_dev_13_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[sleep] ),
    .\dev_13_req_o_dev_13_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[debug] ),
    .\dev_14_req_o_dev_14_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[addr] ),
    .\dev_14_req_o_dev_14_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[data] ),
    .\dev_14_req_o_dev_14_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[ben] ),
    .\dev_14_req_o_dev_14_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[stb] ),
    .\dev_14_req_o_dev_14_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[rw] ),
    .\dev_14_req_o_dev_14_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[src] ),
    .\dev_14_req_o_dev_14_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[priv] ),
    .\dev_14_req_o_dev_14_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[amo] ),
    .\dev_14_req_o_dev_14_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[amoop] ),
    .\dev_14_req_o_dev_14_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[fence] ),
    .\dev_14_req_o_dev_14_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[sleep] ),
    .\dev_14_req_o_dev_14_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[debug] ),
    .\dev_15_req_o_dev_15_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[addr] ),
    .\dev_15_req_o_dev_15_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[data] ),
    .\dev_15_req_o_dev_15_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[ben] ),
    .\dev_15_req_o_dev_15_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[stb] ),
    .\dev_15_req_o_dev_15_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[rw] ),
    .\dev_15_req_o_dev_15_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[src] ),
    .\dev_15_req_o_dev_15_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[priv] ),
    .\dev_15_req_o_dev_15_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[amo] ),
    .\dev_15_req_o_dev_15_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[amoop] ),
    .\dev_15_req_o_dev_15_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[fence] ),
    .\dev_15_req_o_dev_15_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[sleep] ),
    .\dev_15_req_o_dev_15_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[debug] ),
    .\dev_16_req_o_dev_16_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[addr] ),
    .\dev_16_req_o_dev_16_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[data] ),
    .\dev_16_req_o_dev_16_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[ben] ),
    .\dev_16_req_o_dev_16_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[stb] ),
    .\dev_16_req_o_dev_16_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[rw] ),
    .\dev_16_req_o_dev_16_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[src] ),
    .\dev_16_req_o_dev_16_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[priv] ),
    .\dev_16_req_o_dev_16_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[amo] ),
    .\dev_16_req_o_dev_16_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[amoop] ),
    .\dev_16_req_o_dev_16_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[fence] ),
    .\dev_16_req_o_dev_16_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[sleep] ),
    .\dev_16_req_o_dev_16_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[debug] ),
    .\dev_17_req_o_dev_17_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[addr] ),
    .\dev_17_req_o_dev_17_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[data] ),
    .\dev_17_req_o_dev_17_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[ben] ),
    .\dev_17_req_o_dev_17_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[stb] ),
    .\dev_17_req_o_dev_17_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[rw] ),
    .\dev_17_req_o_dev_17_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[src] ),
    .\dev_17_req_o_dev_17_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[priv] ),
    .\dev_17_req_o_dev_17_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[amo] ),
    .\dev_17_req_o_dev_17_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[amoop] ),
    .\dev_17_req_o_dev_17_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[fence] ),
    .\dev_17_req_o_dev_17_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[sleep] ),
    .\dev_17_req_o_dev_17_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[debug] ),
    .\dev_18_req_o_dev_18_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[addr] ),
    .\dev_18_req_o_dev_18_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[data] ),
    .\dev_18_req_o_dev_18_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[ben] ),
    .\dev_18_req_o_dev_18_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[stb] ),
    .\dev_18_req_o_dev_18_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[rw] ),
    .\dev_18_req_o_dev_18_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[src] ),
    .\dev_18_req_o_dev_18_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[priv] ),
    .\dev_18_req_o_dev_18_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[amo] ),
    .\dev_18_req_o_dev_18_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[amoop] ),
    .\dev_18_req_o_dev_18_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[fence] ),
    .\dev_18_req_o_dev_18_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[sleep] ),
    .\dev_18_req_o_dev_18_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[debug] ),
    .\dev_19_req_o_dev_19_req_o[addr] (),
    .\dev_19_req_o_dev_19_req_o[data] (),
    .\dev_19_req_o_dev_19_req_o[ben] (),
    .\dev_19_req_o_dev_19_req_o[stb] (),
    .\dev_19_req_o_dev_19_req_o[rw] (),
    .\dev_19_req_o_dev_19_req_o[src] (),
    .\dev_19_req_o_dev_19_req_o[priv] (),
    .\dev_19_req_o_dev_19_req_o[amo] (),
    .\dev_19_req_o_dev_19_req_o[amoop] (),
    .\dev_19_req_o_dev_19_req_o[fence] (),
    .\dev_19_req_o_dev_19_req_o[sleep] (),
    .\dev_19_req_o_dev_19_req_o[debug] (),
    .\dev_20_req_o_dev_20_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[addr] ),
    .\dev_20_req_o_dev_20_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[data] ),
    .\dev_20_req_o_dev_20_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[ben] ),
    .\dev_20_req_o_dev_20_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[stb] ),
    .\dev_20_req_o_dev_20_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[rw] ),
    .\dev_20_req_o_dev_20_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[src] ),
    .\dev_20_req_o_dev_20_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[priv] ),
    .\dev_20_req_o_dev_20_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[amo] ),
    .\dev_20_req_o_dev_20_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[amoop] ),
    .\dev_20_req_o_dev_20_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[fence] ),
    .\dev_20_req_o_dev_20_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[sleep] ),
    .\dev_20_req_o_dev_20_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[debug] ),
    .\dev_21_req_o_dev_21_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[addr] ),
    .\dev_21_req_o_dev_21_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[data] ),
    .\dev_21_req_o_dev_21_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[ben] ),
    .\dev_21_req_o_dev_21_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[stb] ),
    .\dev_21_req_o_dev_21_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[rw] ),
    .\dev_21_req_o_dev_21_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[src] ),
    .\dev_21_req_o_dev_21_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[priv] ),
    .\dev_21_req_o_dev_21_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[amo] ),
    .\dev_21_req_o_dev_21_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[amoop] ),
    .\dev_21_req_o_dev_21_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[fence] ),
    .\dev_21_req_o_dev_21_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[sleep] ),
    .\dev_21_req_o_dev_21_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[debug] ),
    .\dev_22_req_o_dev_22_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[addr] ),
    .\dev_22_req_o_dev_22_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[data] ),
    .\dev_22_req_o_dev_22_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[ben] ),
    .\dev_22_req_o_dev_22_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[stb] ),
    .\dev_22_req_o_dev_22_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[rw] ),
    .\dev_22_req_o_dev_22_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[src] ),
    .\dev_22_req_o_dev_22_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[priv] ),
    .\dev_22_req_o_dev_22_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[amo] ),
    .\dev_22_req_o_dev_22_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[amoop] ),
    .\dev_22_req_o_dev_22_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[fence] ),
    .\dev_22_req_o_dev_22_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[sleep] ),
    .\dev_22_req_o_dev_22_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[debug] ),
    .\dev_23_req_o_dev_23_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[addr] ),
    .\dev_23_req_o_dev_23_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[data] ),
    .\dev_23_req_o_dev_23_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[ben] ),
    .\dev_23_req_o_dev_23_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[stb] ),
    .\dev_23_req_o_dev_23_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[rw] ),
    .\dev_23_req_o_dev_23_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[src] ),
    .\dev_23_req_o_dev_23_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[priv] ),
    .\dev_23_req_o_dev_23_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[amo] ),
    .\dev_23_req_o_dev_23_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[amoop] ),
    .\dev_23_req_o_dev_23_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[fence] ),
    .\dev_23_req_o_dev_23_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[sleep] ),
    .\dev_23_req_o_dev_23_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[debug] ),
    .\dev_24_req_o_dev_24_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[addr] ),
    .\dev_24_req_o_dev_24_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[data] ),
    .\dev_24_req_o_dev_24_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[ben] ),
    .\dev_24_req_o_dev_24_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[stb] ),
    .\dev_24_req_o_dev_24_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[rw] ),
    .\dev_24_req_o_dev_24_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[src] ),
    .\dev_24_req_o_dev_24_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[priv] ),
    .\dev_24_req_o_dev_24_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[amo] ),
    .\dev_24_req_o_dev_24_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[amoop] ),
    .\dev_24_req_o_dev_24_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[fence] ),
    .\dev_24_req_o_dev_24_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[sleep] ),
    .\dev_24_req_o_dev_24_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[debug] ),
    .\dev_25_req_o_dev_25_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[addr] ),
    .\dev_25_req_o_dev_25_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[data] ),
    .\dev_25_req_o_dev_25_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[ben] ),
    .\dev_25_req_o_dev_25_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[stb] ),
    .\dev_25_req_o_dev_25_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[rw] ),
    .\dev_25_req_o_dev_25_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[src] ),
    .\dev_25_req_o_dev_25_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[priv] ),
    .\dev_25_req_o_dev_25_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[amo] ),
    .\dev_25_req_o_dev_25_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[amoop] ),
    .\dev_25_req_o_dev_25_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[fence] ),
    .\dev_25_req_o_dev_25_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[sleep] ),
    .\dev_25_req_o_dev_25_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[debug] ),
    .\dev_26_req_o_dev_26_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[addr] ),
    .\dev_26_req_o_dev_26_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[data] ),
    .\dev_26_req_o_dev_26_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[ben] ),
    .\dev_26_req_o_dev_26_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[stb] ),
    .\dev_26_req_o_dev_26_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[rw] ),
    .\dev_26_req_o_dev_26_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[src] ),
    .\dev_26_req_o_dev_26_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[priv] ),
    .\dev_26_req_o_dev_26_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[amo] ),
    .\dev_26_req_o_dev_26_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[amoop] ),
    .\dev_26_req_o_dev_26_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[fence] ),
    .\dev_26_req_o_dev_26_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[sleep] ),
    .\dev_26_req_o_dev_26_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[debug] ),
    .\dev_27_req_o_dev_27_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[addr] ),
    .\dev_27_req_o_dev_27_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[data] ),
    .\dev_27_req_o_dev_27_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[ben] ),
    .\dev_27_req_o_dev_27_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[stb] ),
    .\dev_27_req_o_dev_27_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[rw] ),
    .\dev_27_req_o_dev_27_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[src] ),
    .\dev_27_req_o_dev_27_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[priv] ),
    .\dev_27_req_o_dev_27_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[amo] ),
    .\dev_27_req_o_dev_27_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[amoop] ),
    .\dev_27_req_o_dev_27_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[fence] ),
    .\dev_27_req_o_dev_27_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[sleep] ),
    .\dev_27_req_o_dev_27_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[debug] ),
    .\dev_28_req_o_dev_28_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[addr] ),
    .\dev_28_req_o_dev_28_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[data] ),
    .\dev_28_req_o_dev_28_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[ben] ),
    .\dev_28_req_o_dev_28_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[stb] ),
    .\dev_28_req_o_dev_28_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[rw] ),
    .\dev_28_req_o_dev_28_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[src] ),
    .\dev_28_req_o_dev_28_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[priv] ),
    .\dev_28_req_o_dev_28_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[amo] ),
    .\dev_28_req_o_dev_28_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[amoop] ),
    .\dev_28_req_o_dev_28_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[fence] ),
    .\dev_28_req_o_dev_28_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[sleep] ),
    .\dev_28_req_o_dev_28_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[debug] ),
    .\dev_29_req_o_dev_29_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[addr] ),
    .\dev_29_req_o_dev_29_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[data] ),
    .\dev_29_req_o_dev_29_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[ben] ),
    .\dev_29_req_o_dev_29_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[stb] ),
    .\dev_29_req_o_dev_29_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[rw] ),
    .\dev_29_req_o_dev_29_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[src] ),
    .\dev_29_req_o_dev_29_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[priv] ),
    .\dev_29_req_o_dev_29_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[amo] ),
    .\dev_29_req_o_dev_29_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[amoop] ),
    .\dev_29_req_o_dev_29_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[fence] ),
    .\dev_29_req_o_dev_29_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[sleep] ),
    .\dev_29_req_o_dev_29_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[debug] ),
    .\dev_30_req_o_dev_30_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[addr] ),
    .\dev_30_req_o_dev_30_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[data] ),
    .\dev_30_req_o_dev_30_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[ben] ),
    .\dev_30_req_o_dev_30_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[stb] ),
    .\dev_30_req_o_dev_30_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[rw] ),
    .\dev_30_req_o_dev_30_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[src] ),
    .\dev_30_req_o_dev_30_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[priv] ),
    .\dev_30_req_o_dev_30_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[amo] ),
    .\dev_30_req_o_dev_30_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[amoop] ),
    .\dev_30_req_o_dev_30_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[fence] ),
    .\dev_30_req_o_dev_30_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[sleep] ),
    .\dev_30_req_o_dev_30_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[debug] ),
    .\dev_31_req_o_dev_31_req_o[addr] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[addr] ),
    .\dev_31_req_o_dev_31_req_o[data] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[data] ),
    .\dev_31_req_o_dev_31_req_o[ben] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[ben] ),
    .\dev_31_req_o_dev_31_req_o[stb] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[stb] ),
    .\dev_31_req_o_dev_31_req_o[rw] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[rw] ),
    .\dev_31_req_o_dev_31_req_o[src] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[src] ),
    .\dev_31_req_o_dev_31_req_o[priv] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[priv] ),
    .\dev_31_req_o_dev_31_req_o[amo] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[amo] ),
    .\dev_31_req_o_dev_31_req_o[amoop] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[amoop] ),
    .\dev_31_req_o_dev_31_req_o[fence] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[fence] ),
    .\dev_31_req_o_dev_31_req_o[sleep] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[sleep] ),
    .\dev_31_req_o_dev_31_req_o[debug] (\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[debug] ));
  assign n444 = io_req[31:0]; // extract
  assign n445 = io_req[63:32]; // extract
  assign n446 = io_req[67:64]; // extract
  assign n447 = io_req[68]; // extract
  assign n448 = io_req[69]; // extract
  assign n449 = io_req[70]; // extract
  assign n450 = io_req[71]; // extract
  assign n451 = io_req[72]; // extract
  assign n452 = io_req[76:73]; // extract
  assign n453 = io_req[77]; // extract
  assign n454 = io_req[78]; // extract
  assign n455 = io_req[79]; // extract
  assign n456 = {\io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[err] , \io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[ack] , \io_system_neorv32_bus_io_switch_inst.main_rsp_o_main_rsp_o[data] };
  assign n458 = {\io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_00_req_o_dev_00_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1067:74  */
  assign n460 = iodev_rsp[747:714]; // extract
  assign n461 = n460[31:0]; // extract
  assign n462 = n460[32]; // extract
  assign n463 = n460[33]; // extract
  assign n465 = n315[31:0]; // extract
  assign n466 = n315[32]; // extract
  assign n467 = n315[33]; // extract
  assign n469 = n315[31:0]; // extract
  assign n470 = n315[32]; // extract
  assign n471 = n315[33]; // extract
  assign n473 = n315[31:0]; // extract
  assign n474 = n315[32]; // extract
  assign n475 = n315[33]; // extract
  assign n477 = n315[31:0]; // extract
  assign n478 = n315[32]; // extract
  assign n479 = n315[33]; // extract
  assign n481 = n315[31:0]; // extract
  assign n482 = n315[32]; // extract
  assign n483 = n315[33]; // extract
  assign n485 = n315[31:0]; // extract
  assign n486 = n315[32]; // extract
  assign n487 = n315[33]; // extract
  assign n489 = n315[31:0]; // extract
  assign n490 = n315[32]; // extract
  assign n491 = n315[33]; // extract
  assign n493 = n315[31:0]; // extract
  assign n494 = n315[32]; // extract
  assign n495 = n315[33]; // extract
  assign n497 = n315[31:0]; // extract
  assign n498 = n315[32]; // extract
  assign n499 = n315[33]; // extract
  assign n500 = {\io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_10_req_o_dev_10_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1077:74  */
  assign n502 = iodev_rsp[33:0]; // extract
  assign n503 = n502[31:0]; // extract
  assign n504 = n502[32]; // extract
  assign n505 = n502[33]; // extract
  assign n506 = {\io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_11_req_o_dev_11_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1078:74  */
  assign n508 = iodev_rsp[67:34]; // extract
  assign n509 = n508[31:0]; // extract
  assign n510 = n508[32]; // extract
  assign n511 = n508[33]; // extract
  assign n512 = {\io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_12_req_o_dev_12_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1079:74  */
  assign n514 = iodev_rsp[101:68]; // extract
  assign n515 = n514[31:0]; // extract
  assign n516 = n514[32]; // extract
  assign n517 = n514[33]; // extract
  assign n518 = {\io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_13_req_o_dev_13_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1080:74  */
  assign n520 = iodev_rsp[135:102]; // extract
  assign n521 = n520[31:0]; // extract
  assign n522 = n520[32]; // extract
  assign n523 = n520[33]; // extract
  assign n524 = {\io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_14_req_o_dev_14_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1081:74  */
  assign n526 = iodev_rsp[169:136]; // extract
  assign n527 = n526[31:0]; // extract
  assign n528 = n526[32]; // extract
  assign n529 = n526[33]; // extract
  assign n530 = {\io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_15_req_o_dev_15_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1082:74  */
  assign n532 = iodev_rsp[203:170]; // extract
  assign n533 = n532[31:0]; // extract
  assign n534 = n532[32]; // extract
  assign n535 = n532[33]; // extract
  assign n536 = {\io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_16_req_o_dev_16_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1083:74  */
  assign n538 = iodev_rsp[237:204]; // extract
  assign n539 = n538[31:0]; // extract
  assign n540 = n538[32]; // extract
  assign n541 = n538[33]; // extract
  assign n542 = {\io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_17_req_o_dev_17_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1084:74  */
  assign n544 = iodev_rsp[271:238]; // extract
  assign n545 = n544[31:0]; // extract
  assign n546 = n544[32]; // extract
  assign n547 = n544[33]; // extract
  assign n548 = {\io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_18_req_o_dev_18_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1085:74  */
  assign n550 = iodev_rsp[305:272]; // extract
  assign n551 = n550[31:0]; // extract
  assign n552 = n550[32]; // extract
  assign n553 = n550[33]; // extract
  assign n555 = n315[31:0]; // extract
  assign n556 = n315[32]; // extract
  assign n557 = n315[33]; // extract
  assign n558 = {\io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_20_req_o_dev_20_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1087:74  */
  assign n560 = iodev_rsp[339:306]; // extract
  assign n561 = n560[31:0]; // extract
  assign n562 = n560[32]; // extract
  assign n563 = n560[33]; // extract
  assign n564 = {\io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_21_req_o_dev_21_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1088:74  */
  assign n566 = iodev_rsp[373:340]; // extract
  assign n567 = n566[31:0]; // extract
  assign n568 = n566[32]; // extract
  assign n569 = n566[33]; // extract
  assign n570 = {\io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_22_req_o_dev_22_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1089:74  */
  assign n572 = iodev_rsp[407:374]; // extract
  assign n573 = n572[31:0]; // extract
  assign n574 = n572[32]; // extract
  assign n575 = n572[33]; // extract
  assign n576 = {\io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_23_req_o_dev_23_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1090:74  */
  assign n578 = iodev_rsp[441:408]; // extract
  assign n579 = n578[31:0]; // extract
  assign n580 = n578[32]; // extract
  assign n581 = n578[33]; // extract
  assign n582 = {\io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_24_req_o_dev_24_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1091:74  */
  assign n584 = iodev_rsp[475:442]; // extract
  assign n585 = n584[31:0]; // extract
  assign n586 = n584[32]; // extract
  assign n587 = n584[33]; // extract
  assign n588 = {\io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_25_req_o_dev_25_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1092:74  */
  assign n590 = iodev_rsp[509:476]; // extract
  assign n591 = n590[31:0]; // extract
  assign n592 = n590[32]; // extract
  assign n593 = n590[33]; // extract
  assign n594 = {\io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_26_req_o_dev_26_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1093:74  */
  assign n596 = iodev_rsp[543:510]; // extract
  assign n597 = n596[31:0]; // extract
  assign n598 = n596[32]; // extract
  assign n599 = n596[33]; // extract
  assign n600 = {\io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_27_req_o_dev_27_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1094:74  */
  assign n602 = iodev_rsp[577:544]; // extract
  assign n603 = n602[31:0]; // extract
  assign n604 = n602[32]; // extract
  assign n605 = n602[33]; // extract
  assign n606 = {\io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_28_req_o_dev_28_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1095:74  */
  assign n608 = iodev_rsp[611:578]; // extract
  assign n609 = n608[31:0]; // extract
  assign n610 = n608[32]; // extract
  assign n611 = n608[33]; // extract
  assign n612 = {\io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_29_req_o_dev_29_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1096:74  */
  assign n614 = iodev_rsp[645:612]; // extract
  assign n615 = n614[31:0]; // extract
  assign n616 = n614[32]; // extract
  assign n617 = n614[33]; // extract
  assign n618 = {\io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_30_req_o_dev_30_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1097:74  */
  assign n620 = iodev_rsp[679:646]; // extract
  assign n621 = n620[31:0]; // extract
  assign n622 = n620[32]; // extract
  assign n623 = n620[33]; // extract
  assign n624 = {\io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[debug] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[sleep] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[fence] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[amoop] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[amo] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[priv] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[src] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[rw] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[stb] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[ben] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[data] , \io_system_neorv32_bus_io_switch_inst.dev_31_req_o_dev_31_req_o[addr] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1098:74  */
  assign n626 = iodev_rsp[713:680]; // extract
  assign n627 = n626[31:0]; // extract
  assign n628 = n626[32]; // extract
  assign n629 = n626[33]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1106:7  */
  neorv32_boot_rom io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n631),
    .\bus_req_i_bus_req_i[data] (n632),
    .\bus_req_i_bus_req_i[ben] (n633),
    .\bus_req_i_bus_req_i[stb] (n634),
    .\bus_req_i_bus_req_i[rw] (n635),
    .\bus_req_i_bus_req_i[src] (n636),
    .\bus_req_i_bus_req_i[priv] (n637),
    .\bus_req_i_bus_req_i[amo] (n638),
    .\bus_req_i_bus_req_i[amoop] (n639),
    .\bus_req_i_bus_req_i[fence] (n640),
    .\bus_req_i_bus_req_i[sleep] (n641),
    .\bus_req_i_bus_req_i[debug] (n642),
    .\bus_rsp_o_bus_rsp_o[data] (\io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[err] ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1110:31  */
  assign n630 = iodev_req[1759:1680]; // extract
  assign n631 = n630[31:0]; // extract
  assign n632 = n630[63:32]; // extract
  assign n633 = n630[67:64]; // extract
  assign n634 = n630[68]; // extract
  assign n635 = n630[69]; // extract
  assign n636 = n630[70]; // extract
  assign n637 = n630[71]; // extract
  assign n638 = n630[72]; // extract
  assign n639 = n630[76:73]; // extract
  assign n640 = n630[77]; // extract
  assign n641 = n630[78]; // extract
  assign n642 = n630[79]; // extract
  assign n643 = {\io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[err] , \io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[ack] , \io_system_neorv32_boot_rom_enabled_neorv32_boot_rom_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1186:7  */
  neorv32_gpio_23 io_system_neorv32_gpio_enabled_neorv32_gpio_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n651),
    .\bus_req_i_bus_req_i[data] (n652),
    .\bus_req_i_bus_req_i[ben] (n653),
    .\bus_req_i_bus_req_i[stb] (n654),
    .\bus_req_i_bus_req_i[rw] (n655),
    .\bus_req_i_bus_req_i[src] (n656),
    .\bus_req_i_bus_req_i[priv] (n657),
    .\bus_req_i_bus_req_i[amo] (n658),
    .\bus_req_i_bus_req_i[amoop] (n659),
    .\bus_req_i_bus_req_i[fence] (n660),
    .\bus_req_i_bus_req_i[sleep] (n661),
    .\bus_req_i_bus_req_i[debug] (n662),
    .gpio_i(gpio_i),
    .\bus_rsp_o_bus_rsp_o[data] (\io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[err] ),
    .gpio_o(\io_system_neorv32_gpio_enabled_neorv32_gpio_inst.gpio_o ),
    .cpu_irq_o(\io_system_neorv32_gpio_enabled_neorv32_gpio_inst.cpu_irq_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1193:31  */
  assign n650 = iodev_req[1439:1360]; // extract
  assign n651 = n650[31:0]; // extract
  assign n652 = n650[63:32]; // extract
  assign n653 = n650[67:64]; // extract
  assign n654 = n650[68]; // extract
  assign n655 = n650[69]; // extract
  assign n656 = n650[70]; // extract
  assign n657 = n650[71]; // extract
  assign n658 = n650[72]; // extract
  assign n659 = n650[76:73]; // extract
  assign n660 = n650[77]; // extract
  assign n661 = n650[78]; // extract
  assign n662 = n650[79]; // extract
  assign n663 = {\io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[err] , \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[ack] , \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1239:7  */
  neorv32_clint_1 io_system_neorv32_clint_enabled_neorv32_clint_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n670),
    .\bus_req_i_bus_req_i[data] (n671),
    .\bus_req_i_bus_req_i[ben] (n672),
    .\bus_req_i_bus_req_i[stb] (n673),
    .\bus_req_i_bus_req_i[rw] (n674),
    .\bus_req_i_bus_req_i[src] (n675),
    .\bus_req_i_bus_req_i[priv] (n676),
    .\bus_req_i_bus_req_i[amo] (n677),
    .\bus_req_i_bus_req_i[amoop] (n678),
    .\bus_req_i_bus_req_i[fence] (n679),
    .\bus_req_i_bus_req_i[sleep] (n680),
    .\bus_req_i_bus_req_i[debug] (n681),
    .\bus_rsp_o_bus_rsp_o[data] (\io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[err] ),
    .time_o(\io_system_neorv32_clint_enabled_neorv32_clint_inst.time_o ),
    .mti_o(mtime_irq),
    .msi_o(msw_irq));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1246:31  */
  assign n669 = iodev_req[799:720]; // extract
  assign n670 = n669[31:0]; // extract
  assign n671 = n669[63:32]; // extract
  assign n672 = n669[67:64]; // extract
  assign n673 = n669[68]; // extract
  assign n674 = n669[69]; // extract
  assign n675 = n669[70]; // extract
  assign n676 = n669[71]; // extract
  assign n677 = n669[72]; // extract
  assign n678 = n669[76:73]; // extract
  assign n679 = n669[77]; // extract
  assign n680 = n669[78]; // extract
  assign n681 = n669[79]; // extract
  assign n682 = {\io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[err] , \io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[ack] , \io_system_neorv32_clint_enabled_neorv32_clint_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1267:7  */
  neorv32_uart_1_1_e012e0243942cad1e54366b73ee6caff9501611d io_system_neorv32_uart0_enabled_neorv32_uart0_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n688),
    .\bus_req_i_bus_req_i[data] (n689),
    .\bus_req_i_bus_req_i[ben] (n690),
    .\bus_req_i_bus_req_i[stb] (n691),
    .\bus_req_i_bus_req_i[rw] (n692),
    .\bus_req_i_bus_req_i[src] (n693),
    .\bus_req_i_bus_req_i[priv] (n694),
    .\bus_req_i_bus_req_i[amo] (n695),
    .\bus_req_i_bus_req_i[amoop] (n696),
    .\bus_req_i_bus_req_i[fence] (n697),
    .\bus_req_i_bus_req_i[sleep] (n698),
    .\bus_req_i_bus_req_i[debug] (n699),
    .clkgen_i(clk_gen),
    .uart_rxd_i(uart0_rxd_i),
    .uart_cts_i(uart0_cts_i),
    .\bus_rsp_o_bus_rsp_o[data] (\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[err] ),
    .clkgen_en_o(\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.clkgen_en_o ),
    .uart_txd_o(\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.uart_txd_o ),
    .uart_rts_o(\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.uart_rts_o ),
    .irq_rx_o(\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.irq_rx_o ),
    .irq_tx_o(\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.irq_tx_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1277:33  */
  assign n687 = iodev_req[879:800]; // extract
  assign n688 = n687[31:0]; // extract
  assign n689 = n687[63:32]; // extract
  assign n690 = n687[67:64]; // extract
  assign n691 = n687[68]; // extract
  assign n692 = n687[69]; // extract
  assign n693 = n687[70]; // extract
  assign n694 = n687[71]; // extract
  assign n695 = n687[72]; // extract
  assign n696 = n687[76:73]; // extract
  assign n697 = n687[77]; // extract
  assign n698 = n687[78]; // extract
  assign n699 = n687[79]; // extract
  assign n700 = {\io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[err] , \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[ack] , \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1343:7  */
  neorv32_spi_1 io_system_neorv32_spi_enabled_neorv32_spi_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n713),
    .\bus_req_i_bus_req_i[data] (n714),
    .\bus_req_i_bus_req_i[ben] (n715),
    .\bus_req_i_bus_req_i[stb] (n716),
    .\bus_req_i_bus_req_i[rw] (n717),
    .\bus_req_i_bus_req_i[src] (n718),
    .\bus_req_i_bus_req_i[priv] (n719),
    .\bus_req_i_bus_req_i[amo] (n720),
    .\bus_req_i_bus_req_i[amoop] (n721),
    .\bus_req_i_bus_req_i[fence] (n722),
    .\bus_req_i_bus_req_i[sleep] (n723),
    .\bus_req_i_bus_req_i[debug] (n724),
    .clkgen_i(clk_gen),
    .spi_dat_i(spi_dat_i),
    .\bus_rsp_o_bus_rsp_o[data] (\io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[err] ),
    .clkgen_en_o(\io_system_neorv32_spi_enabled_neorv32_spi_inst.clkgen_en_o ),
    .spi_clk_o(\io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_clk_o ),
    .spi_dat_o(\io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_dat_o ),
    .spi_csn_o(\io_system_neorv32_spi_enabled_neorv32_spi_inst.spi_csn_o ),
    .irq_o(\io_system_neorv32_spi_enabled_neorv32_spi_inst.irq_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1350:33  */
  assign n712 = iodev_req[1119:1040]; // extract
  assign n713 = n712[31:0]; // extract
  assign n714 = n712[63:32]; // extract
  assign n715 = n712[67:64]; // extract
  assign n716 = n712[68]; // extract
  assign n717 = n712[69]; // extract
  assign n718 = n712[70]; // extract
  assign n719 = n712[71]; // extract
  assign n720 = n712[72]; // extract
  assign n721 = n712[76:73]; // extract
  assign n722 = n712[77]; // extract
  assign n723 = n712[78]; // extract
  assign n724 = n712[79]; // extract
  assign n725 = {\io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[err] , \io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[ack] , \io_system_neorv32_spi_enabled_neorv32_spi_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1377:7  */
  neorv32_twi_1 io_system_neorv32_twi_enabled_neorv32_twi_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n733),
    .\bus_req_i_bus_req_i[data] (n734),
    .\bus_req_i_bus_req_i[ben] (n735),
    .\bus_req_i_bus_req_i[stb] (n736),
    .\bus_req_i_bus_req_i[rw] (n737),
    .\bus_req_i_bus_req_i[src] (n738),
    .\bus_req_i_bus_req_i[priv] (n739),
    .\bus_req_i_bus_req_i[amo] (n740),
    .\bus_req_i_bus_req_i[amoop] (n741),
    .\bus_req_i_bus_req_i[fence] (n742),
    .\bus_req_i_bus_req_i[sleep] (n743),
    .\bus_req_i_bus_req_i[debug] (n744),
    .clkgen_i(clk_gen),
    .twi_sda_i(twi_sda_i),
    .twi_scl_i(twi_scl_i),
    .\bus_rsp_o_bus_rsp_o[data] (\io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[err] ),
    .clkgen_en_o(\io_system_neorv32_twi_enabled_neorv32_twi_inst.clkgen_en_o ),
    .twi_sda_o(\io_system_neorv32_twi_enabled_neorv32_twi_inst.twi_sda_o ),
    .twi_scl_o(\io_system_neorv32_twi_enabled_neorv32_twi_inst.twi_scl_o ),
    .irq_o(\io_system_neorv32_twi_enabled_neorv32_twi_inst.irq_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1384:33  */
  assign n732 = iodev_req[1199:1120]; // extract
  assign n733 = n732[31:0]; // extract
  assign n734 = n732[63:32]; // extract
  assign n735 = n732[67:64]; // extract
  assign n736 = n732[68]; // extract
  assign n737 = n732[69]; // extract
  assign n738 = n732[70]; // extract
  assign n739 = n732[71]; // extract
  assign n740 = n732[72]; // extract
  assign n741 = n732[76:73]; // extract
  assign n742 = n732[77]; // extract
  assign n743 = n732[78]; // extract
  assign n744 = n732[79]; // extract
  assign n745 = {\io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[err] , \io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[ack] , \io_system_neorv32_twi_enabled_neorv32_twi_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1443:7  */
  neorv32_pwm_2 io_system_neorv32_pwm_enabled_neorv32_pwm_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n756),
    .\bus_req_i_bus_req_i[data] (n757),
    .\bus_req_i_bus_req_i[ben] (n758),
    .\bus_req_i_bus_req_i[stb] (n759),
    .\bus_req_i_bus_req_i[rw] (n760),
    .\bus_req_i_bus_req_i[src] (n761),
    .\bus_req_i_bus_req_i[priv] (n762),
    .\bus_req_i_bus_req_i[amo] (n763),
    .\bus_req_i_bus_req_i[amoop] (n764),
    .\bus_req_i_bus_req_i[fence] (n765),
    .\bus_req_i_bus_req_i[sleep] (n766),
    .\bus_req_i_bus_req_i[debug] (n767),
    .clkgen_i(clk_gen),
    .\bus_rsp_o_bus_rsp_o[data] (\io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[err] ),
    .clkgen_en_o(\io_system_neorv32_pwm_enabled_neorv32_pwm_inst.clkgen_en_o ),
    .pwm_o(\io_system_neorv32_pwm_enabled_neorv32_pwm_inst.pwm_o ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1450:33  */
  assign n755 = iodev_req[559:480]; // extract
  assign n756 = n755[31:0]; // extract
  assign n757 = n755[63:32]; // extract
  assign n758 = n755[67:64]; // extract
  assign n759 = n755[68]; // extract
  assign n760 = n755[69]; // extract
  assign n761 = n755[70]; // extract
  assign n762 = n755[71]; // extract
  assign n763 = n755[72]; // extract
  assign n764 = n755[76:73]; // extract
  assign n765 = n755[77]; // extract
  assign n766 = n755[78]; // extract
  assign n767 = n755[79]; // extract
  assign n768 = {\io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[err] , \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[ack] , \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1636:7  */
  neorv32_sysinfo_1_98304000_0_16384_16384_4_64_4_64_64_32_16_64_9e7924eaddd34398644d20f54977ca62b4d530f0 io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_sys),
    .\bus_req_i_bus_req_i[addr] (n788),
    .\bus_req_i_bus_req_i[data] (n789),
    .\bus_req_i_bus_req_i[ben] (n790),
    .\bus_req_i_bus_req_i[stb] (n791),
    .\bus_req_i_bus_req_i[rw] (n792),
    .\bus_req_i_bus_req_i[src] (n793),
    .\bus_req_i_bus_req_i[priv] (n794),
    .\bus_req_i_bus_req_i[amo] (n795),
    .\bus_req_i_bus_req_i[amoop] (n796),
    .\bus_req_i_bus_req_i[fence] (n797),
    .\bus_req_i_bus_req_i[sleep] (n798),
    .\bus_req_i_bus_req_i[debug] (n799),
    .\bus_rsp_o_bus_rsp_o[data] (\io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[err] ));
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1685:31  */
  assign n787 = iodev_req[1599:1520]; // extract
  assign n788 = n787[31:0]; // extract
  assign n789 = n787[63:32]; // extract
  assign n790 = n787[67:64]; // extract
  assign n791 = n787[68]; // extract
  assign n792 = n787[69]; // extract
  assign n793 = n787[70]; // extract
  assign n794 = n787[71]; // extract
  assign n795 = n787[72]; // extract
  assign n796 = n787[76:73]; // extract
  assign n797 = n787[77]; // extract
  assign n798 = n787[78]; // extract
  assign n799 = n787[79]; // extract
  assign n800 = {\io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[err] , \io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[ack] , \io_system_neorv32_sysinfo_enabled_neorv32_sysinfo_inst.bus_rsp_o_bus_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1708:5  */
  neorv32_debug_dtm_46d1c9a201904415cbd5c7cc672d1649ed497f22 neorv32_ocd_enabled_neorv32_debug_dtm_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_ext),
    .jtag_tck_i(jtag_tck_i),
    .jtag_tdi_i(jtag_tdi_i),
    .jtag_tms_i(jtag_tms_i),
    .\dmi_rsp_i_dmi_rsp_i[data] (n805),
    .\dmi_rsp_i_dmi_rsp_i[ack] (n806),
    .jtagspi_sdi_i(jtagspi_sdi_i),
    .jtag_tdo_o(\neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtag_tdo_o ),
    .\dmi_req_o_dmi_req_o[addr] (\neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[addr] ),
    .\dmi_req_o_dmi_req_o[op] (\neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[op] ),
    .\dmi_req_o_dmi_req_o[data] (\neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[data] ),
    .jtagspi_sck_o(\neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_sck_o ),
    .jtagspi_sdo_o(\neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_sdo_o ),
    .jtagspi_csn_o(\neorv32_ocd_enabled_neorv32_debug_dtm_inst.jtagspi_csn_o ));
  assign n803 = {\neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[data] , \neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[op] , \neorv32_ocd_enabled_neorv32_debug_dtm_inst.dmi_req_o_dmi_req_o[addr] };
  assign n805 = dmi_rsp[31:0]; // extract
  assign n806 = dmi_rsp[32]; // extract
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1731:5  */
  neorv32_debug_dm_1_5ba93c9db0cff93f52b521d7420e43f6eda2784f neorv32_ocd_enabled_neorv32_debug_dm_inst (
    .clk_i(clk_i),
    .rstn_i(rstn_ext),
    .\dmi_req_i_dmi_req_i[addr] (n810),
    .\dmi_req_i_dmi_req_i[op] (n811),
    .\dmi_req_i_dmi_req_i[data] (n812),
    .\bus_req_i_bus_req_i[addr] (n816),
    .\bus_req_i_bus_req_i[data] (n817),
    .\bus_req_i_bus_req_i[ben] (n818),
    .\bus_req_i_bus_req_i[stb] (n819),
    .\bus_req_i_bus_req_i[rw] (n820),
    .\bus_req_i_bus_req_i[src] (n821),
    .\bus_req_i_bus_req_i[priv] (n822),
    .\bus_req_i_bus_req_i[amo] (n823),
    .\bus_req_i_bus_req_i[amoop] (n824),
    .\bus_req_i_bus_req_i[fence] (n825),
    .\bus_req_i_bus_req_i[sleep] (n826),
    .\bus_req_i_bus_req_i[debug] (n827),
    .\dmi_rsp_o_dmi_rsp_o[data] (\neorv32_ocd_enabled_neorv32_debug_dm_inst.dmi_rsp_o_dmi_rsp_o[data] ),
    .\dmi_rsp_o_dmi_rsp_o[ack] (\neorv32_ocd_enabled_neorv32_debug_dm_inst.dmi_rsp_o_dmi_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[data] (\neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[data] ),
    .\bus_rsp_o_bus_rsp_o[ack] (\neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[ack] ),
    .\bus_rsp_o_bus_rsp_o[err] (\neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[err] ),
    .ndmrstn_o(dci_ndmrstn),
    .halt_req_o(dci_haltreq));
  assign n810 = dmi_req[6:0]; // extract
  assign n811 = dmi_req[8:7]; // extract
  assign n812 = dmi_req[40:9]; // extract
  assign n813 = {\neorv32_ocd_enabled_neorv32_debug_dm_inst.dmi_rsp_o_dmi_rsp_o[ack] , \neorv32_ocd_enabled_neorv32_debug_dm_inst.dmi_rsp_o_dmi_rsp_o[data] };
  /* ../../ext/neorv32/rtl/core/neorv32_top.vhd:1741:30  */
  assign n815 = iodev_req[1679:1600]; // extract
  assign n816 = n815[31:0]; // extract
  assign n817 = n815[63:32]; // extract
  assign n818 = n815[67:64]; // extract
  assign n819 = n815[68]; // extract
  assign n820 = n815[69]; // extract
  assign n821 = n815[70]; // extract
  assign n822 = n815[71]; // extract
  assign n823 = n815[72]; // extract
  assign n824 = n815[76:73]; // extract
  assign n825 = n815[77]; // extract
  assign n826 = n815[78]; // extract
  assign n827 = n815[79]; // extract
  assign n828 = {\neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[err] , \neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[ack] , \neorv32_ocd_enabled_neorv32_debug_dm_inst.bus_rsp_o_bus_rsp_o[data] };
  assign n832 = {1'b0, \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.clkgen_en_o , 1'b0, \io_system_neorv32_spi_enabled_neorv32_spi_inst.clkgen_en_o , \io_system_neorv32_twi_enabled_neorv32_twi_inst.clkgen_en_o , 1'b0, \io_system_neorv32_pwm_enabled_neorv32_pwm_inst.clkgen_en_o , 1'b0, 1'b0, 1'b0, \memory_system_neorv32_xip_enabled_neorv32_xip_inst.clkgen_en_o , 1'b0};
  assign n835 = {n458, n624, n618, n612, n606, n600, n594, n588, n582, n576, n570, n564, n558, n548, n542, n536, n530, n524, n518, n512, n506, n500};
  assign n836 = {n643, n828, n800, 34'b0000000000000000000000000000000000, n663, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, n745, n725, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, n700, n682, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, n768, n384, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000, 34'b0000000000000000000000000000000000};
  assign n837 = {1'b0, \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.irq_rx_o , \io_system_neorv32_uart0_enabled_neorv32_uart0_inst.irq_tx_o , 1'b0, 1'b0, \io_system_neorv32_spi_enabled_neorv32_spi_inst.irq_o , 1'b0, \io_system_neorv32_twi_enabled_neorv32_twi_inst.irq_o , 1'b0, 1'b0, \io_system_neorv32_gpio_enabled_neorv32_gpio_inst.cpu_irq_o , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
  assign n838 = {n263, n262, n261, n260, n259, n258, n257, n256, n255, n254, n253, n252, n251, n250, n249, n248};
endmodule

module neorv32_wrap
  (input  clk_i,
   input  rstn_i,
   input  jtag_tck_i,
   input  jtag_tdi_i,
   input  jtag_tms_i,
   input  [31:0] wb_dat_i,
   input  wb_ack_i,
   input  xip_sdi_i,
   input  [31:0] gpio_i,
   input  uart0_rxd_i,
   input  spi_sdi_i,
   input  twi_sda_i,
   input  twi_scl_i,
   output jtag_tdo_o,
   output [31:0] wb_adr_o,
   output [31:0] wb_dat_o,
   output wb_we_o,
   output [3:0] wb_sel_o,
   output wb_stb_o,
   output wb_cyc_o,
   output xip_csn_o,
   output xip_clk_o,
   output xip_sdo_o,
   output [31:0] gpio_o,
   output uart0_txd_o,
   output spi_sck_o,
   output spi_sdo_o,
   output [7:0] spi_csn_o,
   output twi_sda_o,
   output twi_scl_o,
   output [15:0] pwm_o);
  wire jtagspi_sck;
  wire jtagspi_sdo;
  wire jtagspi_csn;
  wire xip_csn;
  wire xip_clk;
  wire xip_sdo;
  wire inst_n20;
  wire inst_n21;
  wire inst_n22;
  wire inst_n23;
  wire [31:0] inst_n24;
  wire [31:0] inst_n25;
  wire inst_n27;
  wire [3:0] inst_n28;
  wire inst_n29;
  wire inst_n30;
  localparam n31 = 1'b0;
  localparam [31:0] n32 = 32'b00000000000000000000000000000000;
  localparam [3:0] n33 = 4'b0000;
  localparam n34 = 1'b0;
  localparam n35 = 1'b0;
  localparam n41 = 1'b0;
  wire inst_n42;
  wire inst_n43;
  wire inst_n44;
  wire [31:0] inst_n45;
  wire inst_n46;
  localparam n48 = 1'b0;
  localparam n50 = 1'bX;
  localparam n52 = 1'b0;
  wire inst_n53;
  wire inst_n54;
  wire [7:0] inst_n55;
  localparam n56 = 1'b0;
  localparam n58 = 1'b0;
  localparam n59 = 1'b1;
  wire inst_n60;
  wire inst_n61;
  localparam n62 = 1'b1;
  localparam n64 = 1'b1;
  localparam n66 = 1'b1;
  wire [15:0] inst_n68;
  localparam [31:0] n69 = 32'b00000000000000000000000000000000;
  localparam n73 = 1'b0;
  localparam n74 = 1'b0;
  localparam n75 = 1'b0;
  wire \inst.rstn_ocd_o ;
  wire \inst.rstn_wdt_o ;
  wire [2:0] \inst.xbus_tag_o ;
  wire \inst.slink_rx_rdy_o ;
  wire [31:0] \inst.slink_tx_dat_o ;
  wire [3:0] \inst.slink_tx_dst_o ;
  wire \inst.slink_tx_val_o ;
  wire \inst.slink_tx_lst_o ;
  wire \inst.uart0_rts_o ;
  wire \inst.uart1_txd_o ;
  wire \inst.uart1_rts_o ;
  wire \inst.sdi_dat_o ;
  wire \inst.twd_sda_o ;
  wire \inst.twd_scl_o ;
  wire \inst.onewire_o ;
  wire [31:0] \inst.cfs_out_o ;
  wire \inst.neoled_o ;
  wire [63:0] \inst.mtime_time_o ;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  assign jtag_tdo_o = inst_n20; //(module output)
  assign wb_adr_o = inst_n24; //(module output)
  assign wb_dat_o = inst_n25; //(module output)
  assign wb_we_o = inst_n27; //(module output)
  assign wb_sel_o = inst_n28; //(module output)
  assign wb_stb_o = inst_n29; //(module output)
  assign wb_cyc_o = inst_n30; //(module output)
  assign xip_csn_o = n136; //(module output)
  assign xip_clk_o = n138; //(module output)
  assign xip_sdo_o = n140; //(module output)
  assign gpio_o = inst_n45; //(module output)
  assign uart0_txd_o = inst_n46; //(module output)
  assign spi_sck_o = inst_n53; //(module output)
  assign spi_sdo_o = inst_n54; //(module output)
  assign spi_csn_o = inst_n55; //(module output)
  assign twi_sda_o = inst_n60; //(module output)
  assign twi_scl_o = inst_n61; //(module output)
  assign pwm_o = inst_n68; //(module output)
  /* ../../src/hdl/neorv32_wrap.vhd:72:12  */
  assign jtagspi_sck = inst_n21; // (signal)
  /* ../../src/hdl/neorv32_wrap.vhd:73:12  */
  assign jtagspi_sdo = inst_n22; // (signal)
  /* ../../src/hdl/neorv32_wrap.vhd:74:12  */
  assign jtagspi_csn = inst_n23; // (signal)
  /* ../../src/hdl/neorv32_wrap.vhd:76:12  */
  assign xip_csn = inst_n42; // (signal)
  /* ../../src/hdl/neorv32_wrap.vhd:77:12  */
  assign xip_clk = inst_n43; // (signal)
  /* ../../src/hdl/neorv32_wrap.vhd:78:12  */
  assign xip_sdo = inst_n44; // (signal)
  /* ../../src/hdl/neorv32_wrap.vhd:81:5  */
  neorv32_top_98304000_0_0_4_1_40_16384_16384_4_64_4_64_255_64_32_16_64_23_1_1_1_1_1_1_1_1_2_1_32_32_1_1_1_1_14ddc86578158058671fcea0fd4647c83d242e3e inst (
    .clk_i(clk_i),
    .rstn_i(rstn_i),
    .jtag_tck_i(jtag_tck_i),
    .jtag_tdi_i(jtag_tdi_i),
    .jtag_tms_i(jtag_tms_i),
    .jtagspi_sdi_i(xip_sdi_i),
    .xbus_dat_i(wb_dat_i),
    .xbus_ack_i(wb_ack_i),
    .xbus_err_i(n31),
    .slink_rx_dat_i(n32),
    .slink_rx_src_i(n33),
    .slink_rx_val_i(n34),
    .slink_rx_lst_i(n35),
    .slink_tx_rdy_i(n41),
    .xip_dat_i(xip_sdi_i),
    .gpio_i(gpio_i),
    .uart0_rxd_i(uart0_rxd_i),
    .uart0_cts_i(n48),
    .uart1_rxd_i(n50),
    .uart1_cts_i(n52),
    .spi_dat_i(spi_sdi_i),
    .sdi_clk_i(n56),
    .sdi_dat_i(n58),
    .sdi_csn_i(n59),
    .twi_sda_i(twi_sda_i),
    .twi_scl_i(twi_scl_i),
    .twd_sda_i(n62),
    .twd_scl_i(n64),
    .onewire_i(n66),
    .cfs_in_i(n69),
    .mtime_irq_i(n73),
    .msw_irq_i(n74),
    .mext_irq_i(n75),
    .rstn_ocd_o(),
    .rstn_wdt_o(),
    .jtag_tdo_o(inst_n20),
    .jtagspi_sck_o(inst_n21),
    .jtagspi_sdo_o(inst_n22),
    .jtagspi_csn_o(inst_n23),
    .xbus_adr_o(inst_n24),
    .xbus_dat_o(inst_n25),
    .xbus_tag_o(),
    .xbus_we_o(inst_n27),
    .xbus_sel_o(inst_n28),
    .xbus_stb_o(inst_n29),
    .xbus_cyc_o(inst_n30),
    .slink_rx_rdy_o(),
    .slink_tx_dat_o(),
    .slink_tx_dst_o(),
    .slink_tx_val_o(),
    .slink_tx_lst_o(),
    .xip_csn_o(inst_n42),
    .xip_clk_o(inst_n43),
    .xip_dat_o(inst_n44),
    .gpio_o(inst_n45),
    .uart0_txd_o(inst_n46),
    .uart0_rts_o(),
    .uart1_txd_o(),
    .uart1_rts_o(),
    .spi_clk_o(inst_n53),
    .spi_dat_o(inst_n54),
    .spi_csn_o(inst_n55),
    .sdi_dat_o(),
    .twi_sda_o(inst_n60),
    .twi_scl_o(inst_n61),
    .twd_sda_o(),
    .twd_scl_o(),
    .onewire_o(),
    .pwm_o(inst_n68),
    .cfs_out_o(),
    .neoled_o(),
    .mtime_time_o());
  /* ../../src/hdl/neorv32_wrap.vhd:195:28  */
  assign n136 = jtagspi_csn & xip_csn;
  /* ../../src/hdl/neorv32_wrap.vhd:196:45  */
  assign n137 = ~jtagspi_csn;
  /* ../../src/hdl/neorv32_wrap.vhd:196:28  */
  assign n138 = n137 ? jtagspi_sck : xip_clk;
  /* ../../src/hdl/neorv32_wrap.vhd:197:45  */
  assign n139 = ~jtagspi_csn;
  /* ../../src/hdl/neorv32_wrap.vhd:197:28  */
  assign n140 = n139 ? jtagspi_sdo : xip_sdo;
endmodule

