`timescale 1ns/1ps

module encoder_sim ();

    // Write your testbench here! 
    


	


endmodule
